PK   u��T��ఒ  �#     cirkitFile.json�Y[s�6�+g�W�]�����CN��t҇���L1� ri&��Z;�1�j1�x�i�����"��� �8�?Ȧ-�
�=>C+�d��p�Ц�bU���Y��<;�y#��^o�JV*3&C!r'�D:�F�	�4w�R̉�,�1�ߟ\�Bx!u��D�A�D���g��c��1C��Œ=-�b9�Q�(Nm$��F2���ǝef���<m!�����B�Q����B�h`�E��dY����e�Xf'���AV�Fs�/.��>��Ȃ�x�Iς��(�#.��]c��]�t]�Y��������!�*��mHT�S�(-C������?��4$친��iH�s9�#Ӑ�q�!Q�'��q�=�9��Ǣ�m�)E*�XGL�dRW�{��d��rf�d�D֘d������df���r��F��Qe�Р[��K>��@��
� ��+`�@�>wE�/���:�Ѿ�vEf[m��eYvc˂{��MH��e	>b74�Z<f,�*lh,�rl��	ߍ۴"۴4��k�;�"�x��[(�9��[� �9�NM�:� ��V�J*P&���[�c�چ!�^W�uC�Y�հk.���z�aUGޑ��-E"K �I�w����~��y�"�)�6E!�DY�I#E�Ժ��>'��h�E�Xbߧ���0�}'�(qh�E	�"�4&�M'��K�+0���AL��
%��K?t��٨B���T���ʶ�)��z#�X�3��Ѓ(;x"!���
- �vU?^W�h�h����z���]�I)�c����ݞ.�J+�-�U��Tu�l>~H���ϙț�P_����5z#�Z�ѽnտx��.aQq�җ3�{�/maP�Js@8'A�`?��y��Ð;Y�3��<	��IU�*ݮ1J�3T�V���CM�}��hZ4i)��z�h����(�s;5��Ȅ?�"����m�l�.�FtGn?�3/tyzC�VuYQ��� A��P�N ���/
���!������:��(���P�a<
�K��d"�q����L�ױ����C�.S�M!�!��`?����Vx|{{�R�����V���<$��u�s�9D;%d~�|,2�҃4�]��n%{��`�r?�`���χ̡��Jf_��覑J=���O8�A�{Y��E����f4[����)������$��d�}�ʨ3�Y5��vJ�4�ߦ�nS��j��zY,��u~�}>mat~߀"�=�}`�P�N�}�2_BF�I�V��Z�.ЫF�Gm_HO	!<���B�\�>����#���ar��T&P�@��aJ�� D'��B�2al��d���r�tC�]G�?���ϡ)�A���tRh��
T`�]��"�|�ߨ���UQ���7�dS�3��~4Z����Gf��qE�_�������|E��PK   ���T�߳�  /   images/6130fba0-ab36-4597-90ea-7b17dabf0cf4.jpgt�T��6���XKq-ťP\����-܂��(��	w�-����\?��s�����wﵲVf���uf�� Od�e hh  ����� ?~���#l���O�����<��}NB����� �� ������91!�rj2R6ZJ��T�/yX^�F{x!.6�S<*B\���D$xԏHp�?}F���9!�3�gԏ�p�$�"ħz���O�����������<:�% ��3��v �%b�Y����h0����@���A�x����n���@�������_�������D@�>��^i*].�Y�N�-��5H~!"�ȝr����˪�.�"��O�PI�2F��7&��_F��~���l׊���K�8U�Z�b-"�X3�#��!v(�©���F��ᔩ�w�W����N�N�<]���S߄�����|`��%s���Ǫ���u��]H���)�bs�l�>���mB������N"i9j��z��QW��*������@��$\p2}��ّiRf�k�"2k՘r������t�g¬��u{cݷ�1��O`�( ��b?�{��y)���J�VP����kP��ߟ8,m�SU���mٴ�p=�P���B?�x����1�+:�R�!��u����k��8���-}�)ة�hI�o�1�������q��hz�F�El��Q�Wv��So�Ǖ|������|<&����1���3�8�9���9ꈨ����O�&Z
O�f���:,�e��r&2n61�^�
�� �,X��������hbUɡ�TZ��bcn��f2T�A61)���2J1���9�_�VFd�
�� �_e�,�fw�VG��@�����^q��X��ꄲ2�y��(�CON�����ŁD�d~�A�F�	��G$�V����&X�Q����0��k�E|���Jq5Z���X��z󿽇]]��d��6
������H�5��[� 6���d�p5�]�1��7Il%Bn�92�_B7v��q�9Tn��,����ѷf4z���b�~lu>i��%��*"���b��:M� ��G�������/�Ot^H._��ޏ���8n�z����qq�!�o��T�����_{�AW��,��}?F��@ގ1C�.�V���V������?���M�����ژG�l���6����e8R^=&�mI7q"a��7�?�90�\K�")^�n���
C�l�� ��ȣ�8[m8�L���9VTM-uU� ��5Է�#�֒���7.ϸWw<uV����<�虝
:�9��Xx������o�4Kҧ�#r2�t��0D��Z`���7���#�	�W@���J.������@��-�ˍyg��f��*�,�`ʜ���/�.�}�ukI�^bV�M��V˻�������j��`���"{���Y>���S!��R:�ؙ� *�U��_X��%���k�I���/�7VT���|@����\)��	�����I�����٭���9������)���K$���o-g���/��_����r�j��^u�I����&�gq���#ƥ��!��\#�`�d��Qq�JZ\�`���Dyf�fʒ�F�z�Z����z�_����*p�9�(#�T��9�����r�YR5�1yaosL&���\��c,�]=f�i�ՕSa^Y���	N�"�d����j'���ozV}c�hXS�*����}o�';s�fw�m"�&7'�}D�]�(b!���{�/��t3�#)�%�>���`	���zA�|�%+���$�lɲ�+�r��F��-��r��T�ю]�#&�bZ_��5�aiwX����-�&
扒�;�gDd�����w.=�|��,Eh�&*�m�h��C�#���wSҭJ��r9�ϩ��U^�M\�vֈ���؄G����o��E�����a9B�7�����R^_��_�xþ�֗v�w��ol����s�|[���k�J�zvHQ�����������=�Hq��m�^��+��nV��9?�qX�V�*���&�2RKvs���l���σ�'OR��r:�����cOvJӮ?�T��U����z�� �р�g����׀�=褐�ˆ�H��Z`��RJ=Q������@��K��J�����}�tBd�}�(����Gc�^��i�٤��s՝?�W[1�?���Lz> s��eB��H˙Nf���Ox]]>0%e�>�*����X��,���;��;=�y?��?����:M;���&@���c{E���f��js/w��!�U��]J�7�.q�S��I^�Ƴ�}����/a8I��i�
����SkR|��ʵ��[/�"�{Cv���N��u���	w<�os�O;�^�p����9w�h��NeT7侊��w��L�eו��C�¤�zo�Ұ#=ab���a��.��{ܜ�;O��@%�*P9ir���h�s�ri��v��Xt�6ػ���]����Xt��|��T�����=�1xo%C�=��%rx��L��d[ui	��ƻ��unj������_��3v��eE��s��?����esY8=���@S�@r�%U�]��M�m�M�h���y|���#=�;����b�:dߦpG�nr�{���P���Ԭ�K!ɿK�?ç�x��D��@_��B�L�[1�5˒"�me�MPm��Y��(J��km�h�7�������x�JH���W�%]���tyW����3.�M���N�D�b��3���_>�o�h�q��������;���� �7����>��j��f�XwNqi �X�Z��*O�v�~T�ڱ��X��:����p��_����.�c�+M���>8�ӝ����������+��(X:�3�m5.d�y쪥����u��Ʃ��ý>�����z0��0��he��Ny��t��U����b��aY��
{�E�/`w�� k`���T�geA4gdN�H�OH���3`��'3�V��S�ֽZ��?i��-H2T�^c5y�?����w�Ϥ���_�b,!rEpD�d�=Q��S�+4wkl�r�{~���֫��g�D^�l���l�-HLJ�b����ҕ�;!-�xYL��� �|ٝ���7�ڌ���8K�@���c,}e�fY]����:��⯊�LM�-�!E㓾K���q�w�p�RpA#]�
�W���Df_�4���ama1�Z_���z�x+����U,T�^� �퓡_G���C�]�4\S�.�W'��1�b���Q
�̵d
�
2E�QT��Ut�`l�"o1��{R1��I�@�����#v���ŵ��`��~XZ�ۍy�����wH��܇���͑gR>┇Q?��:���A9i�{*\i���|�\��U�	�q����MP�L��z6��)5auH{P_����aYEU�d��/?)��0>�@]_|�j����SO������E��U����cj��f�z��.ׁ
=��)\:�1g�x�.l;e�~j�E�<�h��s�-���������=8��������׳v��{T�P]�m���t��JpqQ����\ǲL_� M!(]�b�1���g�^���/�m��&��D��t�jMb�M�"?x<hS;�6V~��9���+]�.�A��rL�%7��r�r���/S�n>�d�.�S�.ͯ����}0�ǊZ�Ϛ	e��u�+�])�Y/��X dc�������?V��#5�o��J���ɉ���O��9�L�u���+a�8�i�;�r���b[��U��M@���ɥ �]���P���X����
Y�����޽�Pބ�/��t� U{*��D�7��c�C��WW�3V
@��N�����_֭Y�6R�,��,��H�k{����s��[������nz&����������t�!��Z�?q�Ńٻ~{D�	밍������I����T~�\�B�ޟj�9��_Դ��S���Ȉ�[(����˩xg��m�XO��M��H����Tb��u�31%��< ~�b�T��*���F�$Ij�����X��o��P��\������@�QX�o��Yu�i�v-i�S��vN�����m��[U�-
vG��҅�fӅ\n�3} &��uN���	S7���x�r@x>����!cw�e>1���Eڞ���f���0΃-
"*����U������8TK5O}�5uxy3�8Eo] �},Ã߄���E��2����Z���5U>4�p��+����������*^�Ǚ�e�,�=k���]'f�Z�>(��%jvLW��)��a�p��o�>@t�s�^W*,En}�5{�&�2��c�9�E���Ǻ�F��Ӫ���E�X�MD�mJ�Aƺ�;�y�~�@o>Z}(�8�jij1(ܢ<VQ�:VrdP��;��:ק��ͿP��� h���M!@�Z�L,_M8Ge��zu�\f�_�z�X5a˱+n�*�>�>�6{��±�*��s��E�rq(���u�n�Nhx�sQ���B�%����M�b����B�٤F�t���N��X���͢+�g�2��/��@�L��xq���V�C��3Վ)�P�>�����(}~y���<��L��:q����r�5���%>�j�X{���o����I@��m����,F* ��aP73Z�T@��슫>��w�x��]�}��۱��6K��t)��eD�o��ݞ�:� VԮ��dr(�}�4��a�N�1�bR�l�u��|�q0��U��Q�0��E�鐫�� _+�M��Bd�ޱ$ܮVl�H;���R�r��ʵ��'닧X�;'���ы�8}��<���~��:j���
��q��y��B��5=M��/�>�T̮���D���/KxW���/B���BH�RSʮWO)�����S�M���"&�Mf�spU��M}��ri�T���j���#%Y��w��hb- ����� -Abo� �W�|�I�0����`{�3��1�;i����������֮���nkԓ��i�@�d�tdTŮW&N<��l����/�v"�gp���#�G�S&t3�w�t) ����a\Q�������� ���i����o$�,� ���V���_�zs����|�?K�����ZK�\�z�CΫb�V����ۀ2�f�LNl�3��ڗaJ%ES|;M�j�i��l�H�U}����!_�}���c��.�z�Į�e��O��4���"�T�ZQ�6��9'��;Ru��D����ɖ���u�O���3�Y��[���gt��0�:dpi��W�%n���"t ]vmQcg>т*"Hٙ;kd��	����X6Q9/��@��^�B�}�����G�}��_�P�$�>�R�6���f�}QYJC���x��C��1��;u'�k�y͞��}:�>i��F;�|�?Ξ�4��Z#G�"[�1:��oT��h� Ro?.OU�����<}g_��$��l�'G�zv_�@o]K��mt���� iA��Thy��lű��w��1� �X��Fa\�]����t����Wu�'K��i��6���;�M�@:�S4j��j}TS�f,�'\�P���U仦B���j�5H�r�)�C�:�3I�I�(�b�0��u�b�	�n:�&��2�����_���EI6���Y<w�s���#��6M���Wy	��O$ޠ�%C�U����<�^��-b3��|����{�w�?B8	.5����J�I� ��K��|��� ��j� �F����\e]3(0s�a�k�W���o�a�Ǩ�j�Ye��h��C�CX���M���4�{���B�E�=�	��מͳ�'^�~/���hy.�-䵣O���_%o�F-���6�EPL�á䏫)����J�Ł����r�r�^�-C�Z�vMM�;�cHH0P-J���h �=<���:P�?و(��V�3�+h1I�� K��R�������K��߇���׿o"���6Q4���]8pKICz�M�#�k�O��&I�.���K�����˹=<��V�XR���1�6bU@e+���T� k�3�T�%����� �����r��(�<5��l���q깂�@qt�T8���L�g���> ��[�KM��,�l�w(`N�
��H7���&3��!6#@i9%a��n���U��`�/��f/ sLy�)w����Hc��}k��9r��h�Hҟ��k�B��
MQ����J�^z6�1B��@O�Kvݣy�x V��|Θ�S�TUH�10N��
�-�_=%�etX��%�cѝ��&bs��=�3FQ\�Ʊ��ݐ���=�����;"��4��]U����w(��`9�Z��:ޓ����V�Rhz���%�`�.U�4�c��D�k�/bI���E�`Ϟˮ�mL��H��+�}������ۮ5*+�.Ӕ���?}ogڽ@��"���E�N���\�o ��;'Q���F��Mh:R�8�e��~��KM��BNQ��|���ה�SrKlWM�A!�!����=g¾Ņ���ǋ��E��Nv=��l���dn�"˯��n
y�� _��kHjG�`��� M-?�E�S�nj�7f�l>٠$���s�ϙt#yt6,�����;Z���%>��S�v�a]���bC*���N��N�g�������i�C���ցxSm�!����Ҵ|�����Dj�o� �Uv/ZR��ϐN�{%��� 5-�x�S^8�0���-��ҔyȲ�"Y/N`Y��6%@�4.�#���)e�"��(�/Id��',ٶ�rQ��k���h[��8�,x�����,E�����{+*��>7�1
����x3�����/C�m"�n�.v���%WxA����D�nq�\6#�ؠʋ�,<���u}uLH���St��1<�Y��o\%���^u��`��!�u��}�8<��y.���&�I@VM�:(XW��8PU���Ww!�c�a�}�&�V|c�}t�z@�Ӛ$A��="�������7�b�y��p;�"�w����?X�f��2y��/�q�qùrubZ�yl�II�nx �>a6�R�{m����Fg��IzьL�F1/T�Ș���6��I�/9q�:�.x8.U
����ޟ�����2�l%���k���*m��(�t��PY�A�FZC�e�W�v�Io������ ��6!�Q�2�w,M�uߗc�-��}7���ja�-���ICF�P�i���p��~_�xZ��V���t��(T���s������<�eA��|����ɻ}G�"`E�����@�chk��>$�tHg|�̾j
J�"ZX�:��Pk�p��!��06�Z�#4M<��k#�
-<��D�� Wc���P�I��c���]��&��~�N���W}��]��AX�BiIH�WO��lh�#�Xn��k��@���햶;@�'~��Iq����l��uVg�H/��y���l}�y�c!�/?��e$D��1��x��}��N=�Z��p�o�iP7��i�VѴ�W:�t�@l�YW0MW��q�z�;��Kv	j[���y��
�BQ��r9�7V����b%6�ߧ�;���S{ǌG������ �dW�HUWOǗ�c9|a�������������V��J�}躨�t,66�����}��j{,��|P���^�}6���J]ؚuF��ؾ0�u���i���ȟt� T0:2�k�**��t'n��p�����"��<�����+) x�����c�O��r.$�&烦��^!&� t�<��u�E����)-O��7�Ҁ���h��o�$k����b1(�t� �R�qه�ڿ{�=���3�y��Q��=5�0͘9Q˔z�|�Y�L����4�c�'�j��a$��=����x��B�ٳ޸��F�����ZEK�EV#H��4�6Ҿ���1�^���P�x(�1��a�����u��y�Ϣ�2��σ[M�]�����ws�����Q�u��إ��g̳I4�pL�і�0�M.O�cc r���}��j�͔A_w_�@��M���B�z�Kl{�qzD�[���b_֤"W���* �Y�&��z]԰SW�\!R����ׯ�/��\:)��1��mvG8z1��{�tf��>4jH�-���ꨢ{hQ�BF��G��>�B2j�c^�H���z��V�8������qǐ�߲T97� J�l�����k���;6��'g���C��<��+1��X9�4��wq���L~��ޕ+ͮyIz`w�����M�]�s؍U���T[�3��`�ya�;F~=��Le��x�2��˭��W�������J��,�?�bF�J̳�N��r
92���^�u}��������}$����t�ёo�+���Jl'�PB�_i� �/� ��ދH��rw���7 ,����m/^C�>qD���@��H�;g1�O��h�k�H���W,G7�����y��\�!��{��Rѝki�UD� ���Ī�X�C�����1!�F_��w�o xh�c7N�'�t[3�f  �x�cG\ֹ��^��+W�><�D�~O�dĉO�9�b�H,.�=�H��/�Q������ގ�}RCn7���S# ��0v��c�Mڼ����ܺ� �P���T�N�¯�_�F0�R�4���T?�O�7���^ &��O~V�$l�/"6�,��'���
)X�I	��U�3������^�zk�p�5��k��~�m����]w��xB#�p<�j�1��������	�D����j����!������e��Ov܍�@�$��E�*���}�|Z�^���o| �ݩ
:�4�d��g�u �G���ޗ��{b�⁁��D'ppn�vg򰖢�:��6}�6ު��h�!�r�Q������������>W�7��"���Vq�V��l�s�i�[��4[wB50�I��~/��9N���L��a��\�U�XH�y_}���tEwy�^{���~
$�G�����,������K�0t�pf���?G��'ʛ�����ߏ������;���Z���ӭ��,(�h:���������5�q���	���a�'
�戃U�"��.5P�M�j����()�/�ٳ�@��Bb�n�	bC�>*I f��Y�!�x�0��4�Wr��F=����Oz 0��A��G��WIʁc�F_���Ss����kJ�<��V/�R��o��a#�aۋ��}}���P{��%��6h��W��q(bc0������v
:]$)#v�eTu�ϵ�C��F�g��o�)]�66�޸a�/�Fݼ hdm����？ʉ����.���ŷ
��Z̝�	�g����@a 9ͬ`�<���u3<�7����WO�ʈ�j� ��n)��X֐��o�:r�y�K���w˫zO6}���
-�}u�d��]�������9
����f�.(2at�}�Ւ��@�����͙��o&Kݿ�q��fo����K�P�b(��#��{��eYl�ϐ��R�[��J�i��{w�饣?�6���TF��3�����;J���vu3,��V�����<]�Y�q�z���Tס����l�U���v��؈�a=ӿ��4~�.��_i����κ]_��D�� ���� ��.�>5;0B����u8T�af-��~��h�+7yA�?_�t� �J#Iq{��	"�<�9����SN�K�R\!���}Pu�k�e/RL@rN����O����>hT��.ڜ�E�B�v罌�ݩ�a��R��w�{"��[����^�Őm���j��>8%��ʮ_����1;�j;�j�8srJ��f5-�:w	 �"J}q~9C�����b2Q���U���1�W�I�~7M��!� ��@�#�F�1Ӱy�|���U�u�7�cz�>�Iꕦ[�4�_��ˢ��Ր��5���E��g� (����T,�lm����M�*?
��Z/Ze������Ǣ;��/-$��sў��n?G�E2|-���d�6Ҽ��.�Q��oSˁ����lLV��4s��v �S �����c��Xt����rr��|���:�7j���L�4\̤�f�5E{�~�E��d-,�������^�t)dF�x3������ʉ��,ӄ�jA�D��V	��p�s����e`6�[4uxP��z�!_�䩑s��Ȋ'�@i<	��x�w�t���u#։2�?�W��J�Ef��T���z�	�`��m=�V�T�c�3����h���X���˲�����B%���Sݧ�u9�D+�������_��m�SG�����Bcǩ,����_}m�'E?�k���:���_Wpk=�Q݂��y���n���
����&�jX�U�;D��n�j�8h!.y�Fm�sQ
�m I����2�X[����� ������7pT�����oKg#S��	�i1�{v("�a|7E^ $�dN�^�4�^x^�%�s�ϖz(z �:UC��,r��v��,�-�K�(���F��o�U��y�]I��p�h?\�nW� Ƽ�g�pE�s�o�6��������T-Z�^�����H�nN�S�m�V��zSZ$�~#:~t�=�B#_J�#�������Ts����C�j��>-��n��4p�%���c��*0]�z/!t.�P�P�4|����k�n�Еd��Z�8�sR���C4�{��]1��$J�o:wG�ҷm;�Ń�t�,7Q?Jm5�����[=Z��r��݅��H^�J��F�_��HZ�� v��t�d@����l�ayJh�����c#���҈w�\�Om��AX��3��<�-�U��
.�����,��.��o�4��;��y�5ӕ��b���s�����Ӛk�k:��j����}���w�nt�yz���\�+;��Bp[��X�L۴���愧�F5� ����!�?_�j �J����,h���+�YH��x��T�~�uD��R�����RŃ0�CMmI 攏�� �H������@�gZ���$+~w�X'd:%�!��BG��[�����~����`O�;����g]hN��5����d�c]s/N��H� s��`;�Y'ba��Y�@ێ`|d����E!'�@+1Hs��84z�D��b{7qRHQk��u	7���ݔ;.p���˕@��)M�xǎ�65����Z"��H�q�}c6A��U��e0ь-0�by�4qɍ�˷���u�?�K���5W�q���J:�EỞ�����@�&�8>�9�9����1��.�/�l��E�g���!�t��	u5<�T�pB���ssh�w-�_
O�Z��O��{�A��gD�:o%�.��$IU��/%:2�y�2�N�_�:`��q�kt��xͰ���܃��B��OǊ��>$��ʸ��`��w j��}V]L�:�[��]���"2J��ۮ�o��X���vߗ�_�@t�}	5dS�/��v�k��~'x66���JnA<��X�P�e�� |��Z�T�wa��D�q�_b�2��j����0��:h��\�OC�����M^�Tl�)�p&z8�����w�^����B�\���K�2�^��p�C����$Xc�s(�fY\��m��Z�h����q�)%k����h�� o�O�����'��Aq�y�\z�{K_OF���Jv�Bs�N� ����N�;O\Tm��L �_�E(�Gw�e�M����-+�yQȈ���+��6�]~'��f���SX㫀���QWהZ��n*�(^���ȹw�օYj=�#��ZP�8��&f�K�Z�}�O��^W��Sf�j��������B��I��c�aS� �;&��]��̂��O�ˆ��.�Dmmu�:Rج�d�:4���Uhkj�^�����#�GE�T�ΨRr�T6���#�_�l��u��7�=Z���:i���O�|X�����Τ��Q?᱁n��)��A}�R�̦8�7T3TT+x�����&����ͨe����A�CFx.�S_H�r����!+��7!�/�t#��]�n�DQjp��S.��/F��"��n�X���B�,��&�'cpK}^=�C��Fqq����<Fo��&}�Z��|Z����5&v��1bñ Rr�RR��:tw�<L�`�74:�Ɉuyܗ���	��I#^��A�Ѹ�3� �}�b�bz:ZrN|�N��$׶Wl,�s_���!]T��u#���5��lT���w l#o	\rP��Đ-O+$����q�HZV�-������i�V�(}�WƮ���_�%��a`q{ِ����\A�͝⣌7��#YR�r}?D{�+?�G���䣡��֠zh�W"�c�6M���eKC�V+��D��&E$?m�>�� �G��݇��3xK�cR/�s�"L`d� �0.�nz�|N��$��A�}��O�\��fFcV��U��d|��O:܃�?�Ђ�C�/>�����ٗ�ڛ�v�N���!U����#��n��G��:��Z5��g�N �H;uڶp^hZQ6�~��=y.3b֛[��G���	!�����F!��.���ڙk������֫j�
�Sm͚�L*H[��Z�� �A��@��A,��].�����Ǚ�t��w$�`�
�J�6���c�'�z���(�T�ˆҍÇ�0�t~��
h�l��l�vA��`�N^8�O "_����&��_�Y'~�q_:��w�.
�t�X�?`���&���EH�����/>�=�D�N��Z��,���m�7���#�E��HO��&R?�})�P�|�� ��a1��M�#�V��ۡ	��;f洇�0?�(W�۝Ң.��`nO�`+��[�+.Ύ��,m1��4��KNb�z��U��s�bԞ�*�~���6k��ZU�c �T`��GJM/X>">!�d)���[*ױ� �SD���&��p�oqV��)Vy�>�|`�� v��Ie\Dd$�ħ��}&�v��*dÄ�4
4����;n|�Ǻf�)mϸ�͓�	�zSVf��/~2AE_��9���zkY��c�eV�#C�G�����K����Zg�vT����ʃ`]=����}�l�fQfQ>;_�1Ao�*�Hp�m���9�0���c��@_zgH��*v������i����	3J�]־'	R�7	+"k��a.��Xc�c�L�������0C�}xφ4�w��qF���~R����-{ە_q�����$�0�l[I��X+�!���P���Oao�ȭ����Ő�^G%����mn������S�8�L��Q}nh�ܳ,����� ���oe-��Ugx/�w�q\�p�dB�g��z�P�.��F!�,��A;�#$���	x����5�r�?N	z�Ƭ�L/�U�0)�*�/�w��s3��v��
�z���?x�K|6.>�*�IK�����w���t��%���ÈiUF-oH߼�Y��F��f��r�e�MvϟE}R����9�p?�`��TB�3(&i�u��$��5�0|�+�~��#��P��%�7�I��Y�6�m{�VQ�t{V����������b��W��DR7N2�L�UQ�(X�{���C���V\��L����A)+Q�<�]N(��(˾�FX���/M�D�9�F��K�W�6Z��G)x}f��pC��.].��)�+F3�*JI�7E�]!ª��v(�XI�MȦ�G!��T:ÂFO�"s���AĖ5��Z������qĥ�����Q�#��o��-��}�c�[���5�K��+�mָ��\t�Є��~�Ck[�ǲ��d�ݺ��� �v�_f�Z7�ova��
h9�̽�4�,`G
}	�y�$P6!�����8Zln�`�ʬ���r:�bm�T��f���?u�l������a���7�C���z�{(vS�K���0=�ﰘd��6��N�-E��x}�,��ɪSO�A�[X��n\��V�c�rW[��@:�y�H�?�>�
~�<�v�m��3�<M*���p�/ܩp��>���ўr5��o���T��P٩�a�*>!��A�!%�]��RY���?�Sy�X�M���&��M��1���s��2<ft�9�J@݃��sW��4E����ZDI�n1_�pn��̒�%�X�"9خ�7�G�MoO
w��VXIH8�8�X-�UYW���>�}���"!_�0TbVEKUҁ�����K���>�9�B=6j�z��O�)�jj���i���r}9(TI]i\iX����[:�$u��Y�_�i�f.(�%�N��Se�+��+��I�\]^)-�}��H�f��ⷈ��3���}|h�-
b�&�m%&!��2�;�lm��H�N@<2Q�$/4������9��2��&���>�H=wu�ѡq�l�4F��S��h��'��s�ԑ�a�(�����!��OAŞD��(��g��i�h�jǱ��Y*�����,t�+'Қm��,��,�sPD�h�<����s��򯬧tQ6�-)"���Ze����g^�+F�2}��Z_ڃ@!���u߮�c�ۖ0���I��LP�w��{/_�\%����������51)�!���%�5�/�:�)\��,Cv��0�R�6�:�l�e�:˶
yE�*g5�����]��m�r�e�B,?�e��7W[s��]�@�h��I%�QMS�w�ŴF�}�z�)c���.{����6����������˔��C��>VZ���m'%������QvWZ�F�/H���,�\!�����߈��r��|J�"�m���Wj�<��px�Գ���ř��}�ef�Ih~ʷ��l�a�S����g�؏�U1�%X~�����r��56�f]x�I���N���^p����k�_h�pE��{gq����d�%}N:A;<m�y�������2H2IQ��3�OڔJ����JW��]�,G[���������d`]���ĩ�s�A.å�D��n��]�9�����6u���.)~�4݄�k��{R��mkwi�
'����:�\�!!�ˌ�7"Z�hˍrѲɐ������b�+���*����mϣ�]^��wCa3*�+�}<p�'�!���LJ��˜�>B��d���%�o�!q[�q��ʲ�XP�����l~��GA��r�t�8Z��.+���xb�g�ѸCˎv���>�Y�)!�1��;`mE�\�Gx��]�|��>�>�&��[��P=���n�c��8а�?��8������Z�S���pl�ہ�,w��K��sED@��n�����gF��ly�u����
n沄�~���%I��3E[�MT�6�S���T�2")t�ԨhsJo:���艹�lڽ�J\��j���e9۽����h�ܛ��n��I�c��(x��P�`��C���Nc+�G�*��M���LB����a5KxO��tO#��|�����ʇI.Ǣ���J�Xfi���򡝺�W�M��݅�o��-�r�����wR�=�?lS�&S��x*��2�vOk��/hPQs\��D�Pcɒ<nZ�QD�HgA~�Z�1��D33��&̒4��������>-��9�[y�8�]P�"F�ֲ���~ѹۼ�2`�0����P���8L;Eû����;��"i����~��	��bl�hV�I�����c�Ґ��S��&�e�J�P7��Y�|Kd���#����1�J�--�b:�Ƨ� ;��&�ۤQQN5k��IC���@ɧb��i9>��;C+rH1�4�Em�G�;m�R��rdϻ�Wq�PL�G������	��y�V�Q����0턁�
�]C�� �����/�Ã�2��ݘ]����MyZJk����[�?8�@�<��*#m���B|Q=Ϫ�	����/�[̲��ȱ���)-?�=`������ݲJ���$�7��>R��i��9`�f�h[�����U�ٱ�N���XY�+cz�Zx���ޜ���4+�<������Cu[�SE�7DB+�7z]/��u=��Ɏ�1hRB8�ч+庙���3��?g^��2���f H
��rZ���ӃeA6��^ٸpt����g�3���ő�ё�NG\���<uD�������"ad�~0���轲I����]y��}߄Po�v���Zɦ�ܩ�.��c����7T9�0��R�{�M�´�L��Wn%4�A�/;�I�q���Q_�����@�VG�4�NR��^���ik��K�q\gF5�,��0��K�H�bd��F+����}���C�כ�u=���.Z.l�wF����V�i7�L���B�8Z`rJ�N�lei%�3<����i��:��20�C�L�1��p�T凰om����W�+�:����ol6{2;>��"4�\[u�r��0�!�b�+�)4�� $�"�+�f�1uk��X��Y�8e�Mu�6L�c)���;�~�!��PA<��X�4�H2��Ú��?؋0���"³�s��IV
��#W�'n޾��j{lW�O�/ŭ��b��W�f]{�"��(�L�nz��+"j9�vߧҷ��?胭R�U5)�z�0�B����r�����+����f1�O���PxR�nH̘���'��i(W�D=���R����^pnR��wn����*���v�=8,�!���Y$��&]܂�ł{ ��kp��������睷���5������sXE��y�Kƀ��Ӓ6k�+��_b���UI���lT8��9�MG,X=����Lk�ަ����ٛ��u%'p�Z�7�0���q��&��.Ng��PZ֛�P�~
�M���V�"��ímPaӺ�P�8�N_��q�ܧgրG�[H׼R8E���F4�>FgM��PjjJ�Α���ڞ��=|? �^y��R\�wJx��2:�g��,{�P7h(j��1�L�����1�˾ 
�M�����/�d�Y�fE�4�3/������\=::�P���cZ��T;���йM����F@�u���_��,h5�c����^i�劷5��֦�\)��U6�ؿ~�D���+���uSp������l��]�<�<f�s5����&c(,��.L��$ߣ,˽����l.�&��3F���v2�i��Z���<p�oK�+�KZ9~Lb�jo��'�Vß�Ɏ�3r���~�	`jz5W^�:����O�m�7���
����"i{�y<�t�,���O�ؚ�mA�wY��^��י�j�fI�%�bX���+e�s���
���3SFۇѣLP�T�&Ȧelį����+��RJ���A�1�$_?q����{��W�օ����v��+3��B��^x�H��z���Ӝ�甧$�G)�">�yP�xɘK�xpoqp{�cM`�1W�DW���~tY�x����t�u0m=�ĭ�@� �����՟(:^�(�)JZn�8��if���>f�]��_c��qY�q��F�J�3��A��mh�W�=�l�C/2P�^R��P�p�T"WT�bN۟i�SI<�t/�rlf ǀk�sɚ���\ӈYR�w��	 `�	6����|f����g�T��K&}�����݊�er��"�h���҈gg�����h���"�*�pl^z��7/���̆SPYM��̋�o>^�����>5i_��@o�r5c�����0���8�(pq���~��qS�E�N}�W�l�IR͑��m=�f-�8��8��ך�hV�T�6u��9���TP�J#⅏If
nj�6cm�#��r
��5{������_C�
!�v�A)�;�|ͣf�6�s�+�s��δ����]�'uo���2�f����m�L�m�xDĲ�d�鑶=X'���l��������e�/̳"�U���{m'���o<�iL��U�d�����9�B��_�SqN��Fݽ�Ȩ�w����[״�V;�z��L-�ϛ�P�YZr+�ZQ��Nzx$0B^�?��5�bKp?m��p}�jeh��<ܣ:�~~_�o�~-���Z��Y����W">>t�IS '��\�G�$��*���c���9`a�B�AH�~��G8�z���G�d�nR�nyE�(�+��7��O�H7�؁t�6N��z3o���j��������G�W�Ɇ/� <�	=k=:(e�f���	��t��ϭ��n�+(-i#��$m{�/kܩcˋq.Ƥ����Y�4t�|�h���`0{��8���	�� !��p��~nq��ӓ��V�ҞE>\��>�`tr��dv]��
��f� ��q���V9 6?�{��?b޽j)���{d��1��*ao�w>�u*�,-]�X���{���$��̙=��}5R�������k��U=x��,��˂>b�S�)��`�zK�Қ�A�4zJS�}2PkV<y��H����b	�ݑ����yQ�]Z�1�����D��}{G�w��w3nE���E�P
=_�SG��B����r��R�Y,(oEݾ��Ɣ��2i���ёe~�� ��b(�U�7}��c{L�57�d7y�lͷ8�e��e/�)�G��1� ��eD�'�fO���Ubk��>xU����4Z��I�;Q�R��η����3�U���;�'ao�WO���/D�a�?�{���q���1'�F��������m��]����������1]\=)�2O�z-��x����ơy+O�(;��/�M�x��~Gɘi�(������ZKHt:�q���� �G������زW�1]o�O�c%�B�����O�����jL��{�C�~f.�Ǆ��%7B���y#�Z�NS<��5�V[%1t�%�ʭ���L�@����� �bZ	��mʽ�Wo ��BNY0v%�E<��k�Nhn��
�5U���+��X�ɶ����,FV1?4��t��OQ�!������ZY��kFm8�� d'� � ��?KMM��h_}�H�O�Qx<qUX��P�H��V��̞ $�@�S�E�*�8���#�;��m��9�!��m>��k=��� ��&����%�lTv[~MY��h4[óc�M���/��̻��b#��M.��FW��G�	�������mC�F�%��ܑ1����}M�)��n��[�ӗm�X�� q_ ]QN>s_ (1A�b���W\ �`�+N�D���g��/�[��K��*�T�]U���`J��4;SE���7�����,�uQ�l!6����E����C�}8��KS%��ý0
z�y߈}� �'�(��ߡ����1�잋Pڢ��]��tg��KSu#<�DM=B�1y��v��G^>� A����whl��� �t겦���L�}��1�槸y���U����e���M�N���%5���J�M1W&�k�������e,�hUn�&��q�=�vr\��g��ͬ�y��^O���&t���W�m��<�k��M��	 J�c���*�J�:�|�:*�Q~�S���.��_9��nۑ��_���\�qm�c���2u��{� �BTpp3����Fu7�oԚ�\#�9�S;9���m��kL6�#I��{�!�ܒYi�.:�5[F$4�����E�� �(������x� q̩҆BJt9�n�5�K�|������TL|���)��,���(��_��(�7s�8jXIO:�&OO���c��[V�_Z{�@9��C4D8�J������W���Z�r�q�&&85ug�{��(��&�VKN�­4�hS� q�зr�C,q�]zKڹ��m�NR|HW={}Top�q���DIi��烼�	H��o��֌д>����yyM�ve��`y�"����JS������;ÖO3�{��K��,��I��C��X��p��+�W�D��h�1+�Vs#�.1�x��x۔k��&�glOuG�\��>1�}"k�dz��`����J�וf������{%m{��!�o�̒ �fmQtz�y|�H������,m��I�Zl��@!2"�]�S������>�b�F�pQ�]�T����x(�����e�F���~�2ՏH�C��g(�B.�;���\&�`����wV�8�j����d�e%!s�n!�����f�Oq-qm��n�&-V��q�B�&������P������40�C�q�Ҭ3���ڨ���yy�d�r�p���C#pB��B��ոu�hf��>�e��p�S0<��g�κ�hF�}R�-�UI�8�y���y'6�k�q�gp��)�P|sEr��xS���2�l)�nx*d�A�=�I��ޑ'Z=�0�Ъ/���&��M��D<dv�[��ӖE協ȿA�k.��N9��O����*�ޥ��d����?:�ҿز��7L�r��b��~�|�isYƯ�7�ͫ1�z��W��T����XX�M��Ua����	C�5�mq��:����'F��$�t@T10t��^�"�rGm��l��_f.PoT�	g%�	�t˥2ݱy��ϥ�Q���(F�᧤�R]�%�Q[�C���͖ �����N�@s�Y������3?�	�<�{G�\	�Jp��O�f�~j{��������^9�!��eb�W|h���Ěѵ�q����v����݀�yIB �[�gG�(�Ԩ�|�bhफ�X�<��k[\%�#"`�zok��dܷ�k�J�1��uʘ�O9�ľ��Ӡ��������H�r�q;���t�)�g
�^sOn�zV�/��,�K64s��W�j#:�����u��UYo��Z����o8/v�ǇTg� ���a�;����5`]g����~�k������߁#��=��V���G�o�����K�!(�YҎt	�H�U8�ؐ���Ł�_�W~�p����,r��*w�7����~���J�� W�����z�IP<5�ČEF��=E�a�x/0�H;���6 J�E�QQ��g��ّ�ȧ�{\̱��\���V�y��t��5�D�t�EW~���,H�#
@��M�.�@��;�7ɬ`�¢���zow�Fh�o�t9��aQ��3s��b�FO��i��Q;��}�;X�b�<1����D�4o�6�Jb���!p¼�h�[(���Z����y�����ͥV<�y��4��gHM2G�<>�ٜ��{�����}�ѹf6M���ǺG ��(?V2���ʵ�Y%���9�'�8=��˯!ML��2�$sS����ǣ����~�c���:��PMa���#���녷8:}�.yG���H�,��X5SB/����9I��z�o�S�M��\��u���1�M�ۘ����o+�C��2�gl\9�e�Ю�χ{�j�3g�d͋QE�_%~dC�:=GԬ� �^�]��d�zj-��u��' ���eo�xh�R;i@_ԙX�"f�b3�mu�A�Nl��R`TO��t��}�� �����1gu�i� �����!�V�Ys�Z�&�V�eh��/쓨��]�|q�Ϗ�Czx��6t��W��A��?VSx��T��������?9. �r�{.�)F�ܵ���F��@vCQɈBd����r����f�N���'��2_���|�R�� �����@�m�I��ܯ���.��#=��O��"�xY�+/�_��S�f���zB!�g�p����A����k氮+��j ��/����|��K�I���Y�U��U��>�d�œņ�"�2�����N����U�a�������:n�<9)�&���֫G��l0�U�$̝�X����Ђ�� yx�~d�}�u�K׫�sÓ暤2�g����fП1�e����f�1=�U����f����*,4�q�m�w���[J̲j���綇�Q�զ] �������	Ɵ�u��&����4w1m����q��(�<_2�yd�lK҈U��[�Rp+֞�d��@}2Ǆ�;�eP��}e��8ȗ�R���� U�Y����K�*oeq�79Z!0��E�W}D,zxl���UX�v2<BD�ڪe�Aj,ǌh���?��ا��@6���P8)�2Z�u��sIzt���-_S��8'��Xi��G1�a�z0��6���g�t)m7b����.;����������R�����j�*6�B�jϕ; �8�_¤�x�\�����w�����g����6�Vm_�-�K(3����`�}	eK�>췿/���$1V�S�m8şL~|g�Z�[�Ja��E�b��Q%�ǹ�x��C�>6yU�e�l���B���9���"�B�)M��p<g��k��M�_s���B�ܲ5E��s��*�����5>�M�ϋh�}��c<%S��������9mHw�FzJ�׼�4𷕪�{��	�\��B�c���ξ��x�*@�>�KʷA���D��EU[c��-x5��b���o��`�\�<�>�;һ�t~�^������58�l`��j.��)�B1�9�f5a��O U��`S�}�<B��Lӟs�^�>�?����_��K�1j�g�e�4��Ȓ�&��q޼Y&�j���O���	��gw6UE�9�h����"���jq���V���+���8�vW�샗�L���!��Y�x�s�=�8���G���eՋ��L�(��A�/��)�e)Ϋ����_�y&�Z�������9�+�x�h������?X�{�������MF����v9Vkx�1rN�YU=e�|V�pO�� GEß6�ԁ�}*/X��>�Bu<���5�'[i�����)���	$:<�)�máZ�`zkw�q�Gj�+�xl��k�87x����j��lH��o�vy���=��6K'��J}�^B]`j���~?X�{*~�p�ֽ�h{�2S�_H���C�D^�LQ��Jm�
��d�υ$�����1���}�A������g��W�oɿ���9�?����6V������N�����P�]�m�M��	����� �|���<��8{Wrɕ��ve+���b!;A��,��!��[d$p�v����jI-!p��߹�� �#fݵ+Qy�(���}^�B�Y���Vʖ�_����G�=H@�,�-���qJ2���b�(�G2�_�h?���}��M��/����㹬Z!����P��R��*h�	8�BcϞ%�P��I��q��g�1~�[�W�E,��w�W~������ID�?����52%�,�42:^��.��/
y�c�sT���Sy��%��(9Ϯ�\��*�Q	�C�;�'��Ҏ��?���T�a���_啟��ln����y��9��q����@e�P�'0�`ԱgP*�YtT���<�cr�yF4;���Ό��kt�<���CW���=��������+wp�X����KO��
���D!���#֮�I��%�>�+�ey��$��.�k��e�~��	�fh��br/r)ڑN��/��\����ؘ^���e���qP�����(a�
	�8R���w"����&��G?�4"����>j��6���9L��>��:)���>e��e�e�fQķ"��Kms�ji����P��Kw)]s��U¤�!��')��yB~�BB��!-#��[�>�I`�v)#\��$C��BxAaY�����n�CN2��Xjj�z����\�hvW��<�*����]���rl�~53ݍS�a)���WC�R�[���P 7���y3{U�!-�<�Ō���]B7�I�_u�tU�?�%���h�Z��x��� �_�����X��S^��a�cb�á�����*�
���ڿ�s�~�
	�P�G�F�E�Zc5�}6Z�n+���W��ګ'�i�u$� R�I<7{�o�:Oӂ	��W+�4Iܭd��9�sY�s��a��Q=��D�8�2��7��n��x��w{đ�`�	S�oQ:�F*�"�v'3�NTQ:,[L�<�bi���_O �7bv3�l�z3�>�U�9����jO� �*b��j�g����|L��!I���K�^3�W�o��`�\���"v)��Ob�||Í	`�cMiN~S����B���hQW�MX7�_Sݷ��+5O�F&���܇���\����\=^�͔�	��k{�l�����|�����#�>�=��S[��h#�n��_2w�pW���D�?�rE�߀�Ř<š���C���xx�Y��F^���2�Ԟ�/�^Q�)�zy��3��^H�N)\*p�O���=�b��'���"C��R���
V�i2�thO5�`��p�U�g��vȮ�&��=f0-,Q�&�\S��y��S.��ϋƉ�+	C�������M9�	=�XM�8O�np�N�#��TJ� �z�NՕ.*����+^�(�Pϼ����\�3��^R8�1�����ܜ�d}�R�ׂ���q���)��% Z��`�9��-�mu<�Y��=��2wd!a��MuNfؔ�)�
i�4��0?0y��'��A3�xx�<���܄���M=9�J������
+[���1�b6s6�쾷	7:���)�wg�3B��ч�ce��2��0T�`*����W�zQ�|j ]0�0
)I�X�֋��#j&�}C���Ј8�+#6 �+G�x�v	��ɂ�>G�ℋY�2����x>

��eOP�U��� ��^�ug�J�{g�i�|x��;�b*H*!��-W`�FW���f&����}���ǻu�7Γ���p��>|6�^)���.-�`\�F@��dp����ױGt��"\�XO �S�ulc��9ˁ��n�#�v��ES<iuCDf�"�0#_]�k�2�)�ʰI�Q��W0�RJW��a�+ǝu����M�Mb������������]�6,�J�_[����<==;d�zP��~�m#X�mx�t�?|��^�r�1#�D7���
g����r��XP/�t[+�*!v��6e�C����vlg�^�B�Sܞɧ[kr6���7�D�:C�ŷ���Hv�J����eM9wZq~�`��R�A?���p�&��������4;c�?��8n��>���}��S["L��u�����KoC��\�LF��U]�<��Y�ֺ���۟�7��<!G<#����)B<����V��IN��W�푓�Z���?hwh|��]����dX��-G�,�|��!䩝n?z�~	�9��%0Py@j�E�D.]z�
���]R��,�C��_��k�|�<�W��-�K�H#wk�!'J��:�q��C�㘾1�!A;���87���pc�~���,�@�H�DXѐ~d��k.Ds[���fFyo�����@����T�e۹)Q�T�uB\^Ĝ�T�.F�5���R��`�
��#�Q�G̢���Jm���iXC\���8�)$C��)B)�̱�|n���J���ǡ�G�W��_R���GT�0y��i�'�KSޯ����R����꙲���~�PAcWi��h���L�r�P��3����M�����������mߓ˙̓���c���g�9�h��cuE0���RE�*���"}����=qr��~~�ٔ��#�|x'�d�bZ5G��|��3֏K���s�h��!KѥW��w'|ݻ!�!|������=h����,\H�g-
_(N}z%�e�����,�'Kٽx7n.�7>�kϲ��SQ1d+Dg�+<����V?�Z�(i�1b��y������t���;E誕6?�@d��Y����>B�G���?+-t�fC>�9�0#�PbE��={��6�i��+�r5<@�U�f���s/&;U�R*�6�C�<�#P(G�;����H���Z<ʢ/0Vx��XzW$�*�:Vòs9��eW�������ԑ���M�ٴ�˿"D�4�V�+�@��̫&\	�Ԋ�>����t������{;�N�����-<�+�W���C<�؉JV�rj*��&�ͭ���f�U��� C�GQ�������o��� ���$59ҹ�$���cìp��ڌ٢ɞ�4C��U�B�<^�І!�����#xF���3������}�P*i���=3e�3�[���}�6�6�UU����=W���޸C��3��*>B��3����"�:�u��1�u�d����!b�p�m�j�q�W��Js�%Z/t;������;�I�0�UXW�;����m��gng�����h��	扁ҸX�����oB�Xк:j���p���Sa�.==´ ,x�,���%9�[AON�/��8�A<���nmHs!QK�{�ʘ�f��D?��~��#\/������Inw6@z��f�zk����x��[~%vs��.H�s�	�^?Z+����P��v�w�>#D�In�TK4ҹx��_��#���(}�����ɋC��,J��������bBV�i����_�(���iO��/Y��x�i�;V��S4����)~���;k���-"�tk�t��p����@����m��K���yi���;O�����k�9V��2�݀��,D-�����C����kяf~�xMg����i��(��ڱ�qGlȿ6�zN���¶�ƙ���)"ֽ2q �͆R�fv�����2/`�����jHEo<!����^H�@��<�s��J��U���yt׫�pXؘ��_V��?��S��P��[�ý,��j�����U��5{p^��b`�?�S����	Ƽ�yt�*�ZY�dƳ9�H_d>FC�M��""��#�H��>��h�jѱp�Ü�YI�����7-����A��w���+�>=�X�S�zw�X1�;*j���
��n�����-�TqAu�1f�0�L]2ٴ~��i(م���O�_"Jt���KE;\�K�P){��Җ�~/��AE%��^i��V���������X�Sˣ�E-n�Qt����B�	��Z��-LG�eS��AL���{���t��
u���	�L�W (Hv m�d�{�n�awJv��XV4v�p�7-�)`�D|'��D�2Pm,�j2��%����� 6���'~F�rF��XMaTJ����=9T�INd�ĭC�{|p�h���"�ħ"��Ӟ�#�њ��HP��/��$i���ܙ/��;W��T�J]���1�ɔb����@w���)N�e�e1�B� :���Amx��F�"�0!JW�����ؒ�)8J!P�{r��f+���'�P
���4���~n�B������Jdˏ�S�F����ڍ�_z�"�0�Z:��Ms�`�L:C��x���!���|j�5��fVK�c�tk���|����w�gls��O l��'@$��� _(a�ٛv�O��u��c#X]��F��9��>���?�1��w3^��i��1�_��w�lj�tH�L�U��������Tʅ3~:~�����8����\ُ��y"C��.���>Ў���?[���h����N/4��
�r�bA�lxm�O<M����|��}Βմ���ã�Ӝ��*�Ԑ��}s��>\��O��,���	���fz�Y�j`G���IY	�iLLzIg�FQ��_*=K����Տ����t��Y�j=UR>@�TNаn$�� (Ĭ��Sl*#2{�nң�S.��A�8W v8�'��EW$���ؖRhe�lō��kj�hgo=p��m!��(��7���^����	a�a��O�5~K��U"uD�nԗ?YŰEg���f1Er]"k���>�!;� L8�Zu5�$�gI��*7$�6=6^ S�3Q�pjA���R�)`�Vf�oԊ�¥*fſD�SNo|ɣ,�Y��b��p�V��i��3<,;bE��˧��p���h%6T	[��7�@�?�K�����vs�W��)�(ym���G%�h�6Ǘ'mQi�LI�1���
��ԾIo2���0Ģjn��%��g��?×��\93�G�E"s�ŶӜ����۶��-)�/=�*i߳A����)o���`AmyaD��J�����z��Ln�_h����Q�AI��Q�zZ�w��c%��y�?���P�����#��
�!"F�Y���ߓ������A��2��%Z�iă@-��Ĺb}�$����H�oy�ۏ�lv,�[2u�����=E�+�H �e���J�[�s���T�إ����?�tY*ODt.������	������(��@���C�M3�%�t�]��j�F;2��=���卅�j[�h�`�G;33�����	�O��y��~��;�?W´�D<�O�.�J@��su
 ����;�٤ΎD��=�-h���{˷���d��s^L�iV���'Â�_����n$*)�&q�[����n�8��_<�C�u��y}.ڭ�^�էM��Ruѡ�r݁�l �V쫏+L�ջ���K�W�rˋ7{H~x�IƗ�0?kV�s�'i�Xtk�⮺�"�]b� ����)��YЩ��|�2����@���_؏\44�/�q�؈��{� *Q,��Xh�u��/��a���m��⧲��[C��i��7���E��ծi���)����I�6ߚ(�KӛN@���tۍ.@(Dʺ��H�Ji�ެ!":3�ԯ�ςݐ�� �ȷw0����	 �����@]�VЋj{�o,U���.Y��?����h,Wy�*q�/̒B���	
��\�.R3&|��>�1�J�-9[���v�U��LXK��e��4P�1�/�zSO̵I��H�fj���ov��� �<�h*7DN��Zi\&�wq'u����<�5�s�s2��$l���[>�����sd�(�ߧ�K���3�����S�Q�����0��Bf'�ҁ��{����#){�7�u�(y<����(�/��r*:=ߌ���{��Ģ��c����mn�����g�ڨOg�����i)쳙�w���R�O�&S��r�Nc��S����NZ���H���oâ<4/Dt��?��{�����Le[���w�?���)��^}F�7��"rF��Fn,���ʽ�d�g�����a�Wj�l����*�0�3)7Ȓ�$��Cv�/0�Ȑ���{���' =왎���ܡE���E피y}� ��'@����}�\�G��6����m{�]�d�Bf5����Cv7��}�F�Fn�k1�7��\ԡ��i/n7�ne?'2��,�X������ Ł�ĳϊ!�g�ϾNg��$�R�Z�-�(��{0��I�ҞN��$',2����ڗ"�g8Z�4Z�*.���A��*��iL.[�[�~�|^��Bx����?��}���{vU���TTL������V����4	Z;��%�����L~���	C}�(j&.GE�VV��1�݀ �V7Y�g��ylv�p	��k���������棿�4�3���J�����d��D)y�@أ��B��1$��s������z4ɷ�=����$�dͪ�SI���4�⎧�̑
d������,���)&��pb�q�ľj�*��z8��$"�[	{5���5�T�va���<�2,�42L3q?ΚN�s��*��R&�ANC�<���$�i-���&�x��ϋ ��.�d|}���uڊ5y�ZF��i�o.�
��������I� �zp��I_���Y���䐅���j"Y�W>;E�ru��A2�|P�,L���J ,�F����f7�@NoX�|�U��A�cI�K���.t�R^$F���g�$�6�tg� K���DfJ~kn阼*.�	H2Μ��_A7UKµԻ�̞~]�ٛ�;�_>�9kfk�F#�_ �lFR?�+��ןK&�/�a3��1�`���K����+�ƿ� �*K���Jcቋ�.E��ԓ#�H;pc��Ш��Ѯ�fi��H�%�� �h�s�g�����t�̓��l�*b�z��G_�a�=*��@����*�Et/;;66�D^�_Fs]�xs����cg�I�s�^��	�-	#���u���w!r�qSՄh^���V`�}�vZHb	LB*�4����D%����G0��`�G�BN�T���>��r�z�J�5�ܥc��=�8��K�����)�İ(\��Q1K8�8���}	�s��r�� �Z�5y 	�x�/P�?n�X:�mƐ��*
-�����VDb`J9�N*�v��@D�`>/��;�Fc�^o.C��`�	�Q�-���C�p��	�U��Hk�S�+�G��7�E�mV���	��97�\��2I����@�R
��S�x���:�����׎m���%�<�xl��1+�i�������^+.pi|)1�&a�\�@�y�\�$��z�f|t�;�)zV�$2�9H��T
"7{� �,�K���Ax?wذ6�7��h���x�i�Oi�]?������ E�j���� �@;ڕ�p�����G���y��ǈ�h�^�yq_��>6|��Fw����J�[��R
���>�D&HY�r��Z������9�uٷ�q��׏W��:��xc�d+������| �癵����FW�ՙ0���Z� �����kN_�'��Uua/��#HL���5�L��s�D����l�v{�J�L\/�J:�L�WI�\�����u�
�I���$!w��\�ω��,=窄������@���Am��yxQ")(.)((AaZ����C�\cK��ZŔ�Hy��2�bs����\<���/��C�VWW�Y6���iدm�]���?�F6�/���	{A?��Y7�4ӳU72�G���*��%�j�ZyT��3a�k�������2Q���_�@:::F��4�b����X\#V��.��3��h����|�EcZ��J�&���㧸���Oh7�V�U+4+r���<���1��v�8R�ƶ���V�[C�+ô|´߷�1i�Ao:�+�Ug�zD�҉�W�<W�w;.j�)�́�֏�>�3?=��-kƯkE��<��DS�ķ�����.�U��4��gR��I����-�D�A��G��Z�8I��T��O������q"J1%%����԰;�D�����T�7��D�=Z��=�iؗ
�zP�3��\QͿj���@)hO#���K��+1��ef��m�`�ڪ�t#p�T�k}��^Q�iP�x���#|��:<.�޽~W-�����]a_�>���M]&b{��Y�u;�����3�)--�^1>;���'���
gz�U~:���8�J-=Q�z��S���Z{����s��t!ł����}��=RS{a��1���a�镖ӻ�b5�|%5�@�3.�h�Ts���`��O~�JBRc�f�������&���������e�@���ĳhj�fB��]��J˖�w���d�-��h����g`nys���-m��zsL.�+���Q{�N�]�!��4@!�.=5:0(8�X�S�A ������u`���-M���l�毋}�3���8�Mc�Saݨ�����C�+�*((&�O�@4䫦N�H1��yG{!٫��Vpa|�x���o������	�ĞG`�� �r��V�ӭ�*��\}� A��x�@NY�5ҫP�	����і�ֳ�f#��5��q��s]��I�Y澽/'ݧ|5�j6���}i�;�Ա��ۦHf��O ��.���g��5;[�'N�������Ѡ촻����K� ��y$0�3��ʞH5/�M��:�1�;X8����Mm�>zSv���$W8C*Bb��u�-�x�O�K���:�I&p��y��N!��|pS&��c�	��<𻠱��	���(V�E�H�K���a�܀�n�-�*tJ]���̙���`A�z��Q�9v���o���2��op�`GI�}9��ۡ��sR���L�}�ʧ�0�'�-��D�AHb��|�XD���H���%듵H[�'@n�^½l�k�2��5=���L���`F�=�Ŧr:�����4��\�M���Ƿj��{I�5��*_��3�F_M���1��hU�7�%%��ڀ����h�jھ�U��7e��Rr�q%��Z[�Ȥ1g_�(���l��[Bn���u&��#F��J̷����"��1�VK�V�0{���Ϸl��m�3S���㇠��>�26#廥����ۤ�����{J��>x��)K)R��{�hg��4���A��+W�X�7|���}�s�ͩ�3v�Pl���.v�/��V
���b}���V�=��� �;8����7�� �Bh�&d�g1N$=+^^�\��8��؂�(��`(��}/c����CJZz��+�G����G�������������)}�
x�@�a��������F�?)�'�c����蚏����u�i�eߕ�m�{仼ȫ�\r�h!�u�Z�|@�U@n�ܹdO�ýg����~�U/%�%�bMak����M2>SU�}���q�5l�W4�C� �-�Ѽ.Rtn:Fa;�����s��Q�	�&��kZ�6�|�e�*{��A����W�����k���Ӧ�����r~4��A�:��[���=��؍]�N����nM�s�L)>r�:l��\4��m�&}�x��f9� {�ntՑ�Z9�y%>*�g��dF)���L{�Gmq�q�R,��h�-)�Y��%2ۂvAJ
G��FѴ�r�#��O��b��<��w�����'��ƾ�"����~�Y+����?��ƥsk��cwg�~q��fa;7�o
�7�T���N��n�ۗ[��\{���7Gi̺3��S�/n����ឨ�*�b�]�=>�XEժ�L2
;�sz���9/
�ӿ��7��hr�&�q�B<�u؃tm96�ex���P��%�*f}D��q)�X;̟�P����T��8��`s�h/ܵ��pYZ�����xl��\�d�g�ӱ�-��y�ʴ��v���B��wd��������(Yv���ʭ�I?v�+X�%�O��_�9h SW@��T���P�l�EJ�����9���M���T�}o�lBq.Jc�Q���)Q��K�Q���ԡ$鉘��.9����BҚ<���
b�!�+!G7d��`��#v���y�^���#{TE|t4�]���q�4�q�w��kFSIԧ�}��f�3�Մq��D|D�9�]Q��b�9��:�75��4�e�hv���֭��� �p0��s��i�������S�?F�M��r�4�v�;�a[�{J�}��=��7�z������]���YJ�c��lHY}�j�a��p��#�8����Ɖ��D��{>y펜�H�(ª�_��{6W#�+O��
�Ǡ�����7,���M�����
�ֺ�)���apw+P|ܥ��[�R���^t��݊��N)
�Я����s�{%y"O���4r_�5�	7I����0����ơkʹ�҈ �|RJ8o����.Io��G/�(��/�|��X����^�^*��R�I�J���F�7}F�6�X�^��ʗS��/ޚIC5��N���XXY~l\}�$ۆ_̕��G`�S7I��Ax�8����!Q�ͬ�������5Fb߄���>}* h]�I^(��I����:wnY+w�=��֙|,x�l1_x�5���w=7��2Y?*)�,��<�K�kؾ�*ט>��U�'dpdi��o���Zd9�lR�P7ʞ�?wwΈ��:v�N8��d�1��<_���`�����,wssL �f��{�up�K����������Qp������'1i��G��|�� ���),��Α�㪔��f�5���� ��s����P�N�_�N6�ߞ�ۜ��6Zs()l�S��+1���3�������Νف�ww��==붿%S��ɲ���J��[�vy	��i?���,}��o��Xk�D�O��d6-� ���ר��r���%Ti�@��o��^Ox����M��sNT�(a���Z��,ޔ���kyv�ۭ3��,ǿ(�g��g���7����lOo����}"=������ܮ�׏%��l�ݶ�\��<t��v���L����l�	������y���F�������?�L������R�� 3	���ޟΛf67x���.��k
��0��j��u��is���rλ7��=t�K�r�-��gCO����AR��s^ ɪ�E��ݪ�%W���Z׿$�����8��BS;"����$?
��<G��?��>�u�͌�6}?��l�ݴ���(�ţ����E�ʨڲ}�L �s��`I<��ų����9�CBDAB��{f�7��|2Z�x��a���K����{W����4���j���������^��9�b=-�����)[Y믟��	�H]Ǳ�]�;�����W���[�A���\�P�FFx���5�1�j-x�v.$�9.*�\��"6�Rc�.�*kK|�j.�^X�4�6�]eo��l'��'�N��c&GQ.S�^C����W%�8:�k�g5�ƙ�������nv��p�6ڈܨ1�1�eg�A��X�L`PmҸ�GO?�KTc�j��� �{} �s����|dJ�-���]t�-�Bʌ�l�䍬_�J�4$4����:�O�i`s��@INb(`�~�s*�/��H�b�p�݁yV_<��)m��p��_���X�|�tb��
��ᰵq|�g���GW�`��,������T�,v5Ԓ��ߘc��`;;�[�PS�M��_���&:�<a�Ý0sC>YxWQ�X��M�h��%$G2K@6L�{��'
­�H�9=���v���8�.BG��{}I������vs�)��%��d�Ճ"��`b@p=GBw1�R��E��pj0Z����X���#��뮝lJ�b��OɵN�����8e+����M��?���8�DBE|��|���@=� �?�=��`]/��(�&�Y����pA�_1%��.��������
*�6@m���8�k��Emğ�j�p�v0n�-p0���y���݈
�!.}����V�SԤy|p�VL��Uũr"�FɃ�1�|�Գ��`���wqW=�����xf�_+�-�y�;O���JAb%���`��.k��:r�i֒���9��B;W��ʔQ_��խ��Y��I���Q�bL+i�5�[��a�<J[ï��!��[�a*+�e�<IW�A��	}�UE�KZ^�߶�1� �FQ5O���Iy�R���1��n��1 �Cǚ�h޲kAa��S�I�j΢N醐e�J����l�}�Cw�$���f���|�'X�ͱ{�f��I_��-_I�+D�w����CD'�Kc�@��7�$!z����N�Kk��w�=(�,1�/�b݋����; ������I-��_��X?�J�1α��������J�c��md�>�y��`cXM�O$�P��!LΚ�¦��������	��y�������H u>GM���cW��/#���$�t;����H]Q�6_%R��#ɂZ'���B��@h��"�(el��*�, ki�hݍ��3
H�g�qX��^I8��#&��% >����e�MZ�A��ü�r~e����"N�~���Q���C�L�������$fHtv�X����#��
91�jƅk��-k�	ʌ3�2���5>⃔����a�Z8xǥe����K�
�(�O%�nѰ�(�f�p�K�.�HqN�oF�1���EXc������K�D0	���1�����RXF�����mR'L�� Z]�[�s:&�'r�\���c	07�^���_e��&�F7+�n 6L�����i��`+��2��&s�3��_�~Uk�p੗�>qJ�F|����EwS#�m�P�GE����h�8��1�r~�=�����c�3���q�j�w]v��Q&B��N�L��1wf�W�����(dlF�4�v��Xk��եw������	7݌	]�Կ�L�tZ�g��a������`�n%�vؙV�c��O��!�!Gz��5:�&�p����0>��v������J̌3�4�������a���-N���ŉ�c�(���.��e;:���KS)��RQd��� ��c������:S�p~e�R�  7�_�x��D���%��� E]����X�UM桋��$Yb3\�fY*|f'~k%4Z�.�e������U�(�%��$*�@((��1b>r'�� ,����'*�m��,R�q)������ܬ���Z���I��b[ۘ��Gq,��S_>�R�5�f��5��$}:���V}jIm	pQ��ށ����nU�jomP�>��+j�h�H�'��-�D�	o��>a�3�����T�,k����)�OTֵ�̲��P� K��[�ʓZ�2�z�؃Ẫ���E�t�'�f��R����0����I�99K|^�yf�u Q��G�I���}'�^�b!'t;$��g����;�7F��9r�a%�h2.�|j��^�I�܂��.���j�E�jx�s{{����E�}cn���}gI�f�m$�(���#=yri)\��r��Gtd����V��%�P�pT���/�-E�%�"�1\Q��0�q�('K������!��'6����Xe��Z"%*��<n���>�K�ɜ�,�dXJ�3�H
�H*�KH�F�rx�O��8&#%��3��4�&����&�ӱ ?�a.yz:�i�i��JD'5�D�@Kl�5�B#�,���}�{��Is�D®��[^Y{ q~44ˊ��z��q��k��mN������%���LU�^�o�?|v�'}^�\a���$�}�b{ɴL焗�l�V<�fZ��Y`^���ix�׿/�R�[�Y~��	�[�&k0�������w\�d����V̆l����֦��,�o���@%�{�ȁ���>ްܜ��HW2�[��]�4F<��+�ΐ�]E ���\�U<��Q� #]���.����r��]��Ye��T+=��x?e�<e��E�I���[ѯ��i�\R����@}b0�9N��FwK5�F�^n���T<|�9¸잷yN��3�Y))�-zʭ�|�t����&h+�����)�ǰWX�������!K��_;���5��� q)�����Tu�6���=�cgL���+_��I����`�$p�����SBY� �k��0�q#�r\P�����n�v�Ҡ�Zb��P�Щ ����N���:o�m?�IPe��?}����y��hL45�B8 <#=���y��Y�-�Sg���8w���a�����cTŚF^f���O4��te�)�"B��_l1Hj���=�5~ݤ��I�u[~�	�(�qHE��@���IgLY?���(��e��ȇ��=\&����o��]��<�%TcnzjFab�d�$�;���$$-��s��"�ߤ�1w�Wk�I��f=K��~ə�����U�q���l�"�=�*�c�0�	�9�		���F�s�vc~���^8�r
[�}=㲥@)cw"t |R�� �"˔��q����sR��.�n�_d���c&�܍\�,q�7G8 ŷ��Hm��k��Pg@��eiNGQ㰸��'�n9�}{�������d�t*N�!���ʱj/�F�;��qZ=kw#4�������Yc���[�dWXޫ�Z�Ű���y�r���0����6�tt�M��[4��cc�h�����[�N�!���D�^���|�^��	.�e�S��x���[| �\�[�O+����d�م�X�i**{'r{���k�����D���*�ĸe���{JUO@����^Z�0��n�ɟ��"�+:bs��L��+�)���[b��^��NM}�b�=�49�u_!|RK�> 4�^�/A|{��/Ě�'#��Pu������_���2P�,�H C��S'}�Q��BvJ�rCwm/��"w1�E��<�w�l��#ݳ������	{`��а�/�ɉv����x%_hݿ��?����?ŨlΉp�����5(}��;W���/��GDM������e���w6Y���z}Wb9�<ا�"d�`��>�i63�K]�C��"��^�ݤ>i���7Hz�;��_ 2�@?��%cb
�3���h�{�~�L�4DX޽m׮h������\x�(�̀�b��q���摐5���`yI�)_c�w:�rzD���<{�xW�We0�b��ĴR^`�a���9���B`�X��L��
�8��[��)��cȃs�B����ƅ�8m���3},�3ȫ^�Qj
|�3V"8;Z�/V���� ���LE��i�{k�:=�QΫ$/�I��_W�51�@_O������@��%H3K���@1���AP�σ[a�⭸Y��ҏ�<��ǜk�c��ٜBJ)a� ����K����l|'9z5.��
3���Bq��"��� ��4��N,:�<���g�a����\�
Mz��s<�`�!���^��"
f�Tq'<V�NJ�E$+��h�����ڣ�;5�H��Ui~G9�c���P(!"U��i��)�dv\ܡ�����Y�T�I����qɔ��)?�'���J:	O��	;%� ��8W���8�@�E�����!ԉ�q��H)����_�B_4u�(%��p����&��ݤ;�xC�T{���1��w4���ڳ�/^L(�K�Ul]V��>��m;���L�*�tKD��3����l?og@��"��/�����t4����������»q�����X|-�W��W�p�fv3�2��]aE����HY����#1b8g�8�<�٤TݰCP�˵��q�Vx��"��)3���� _1��O�g�@�v�<�X�k��͗�<��%#.�!G2YI�^�.I��æ>���?��{�b��8L�k��~^���Yh���U;[��M,VF��b�$��x.�O���K�nyXX��}��b�g�x��̄x�S-[��D�E	\�F74���
�1"�R ���<�(����������E/����������1k�������e�42�3��gW�_�D����\r�r�c�?'��E�I{�Ӆ48�i'|�pE��q�&]
A�*1.ϑ��NM��jzcy6N7��in����$&�	�m�E.Uj����C����F����
l�ժ�,oc.��g2�N�P6KmE������^�*	f������V��0, �ܢ]�0�<�����
��`<F9�Xe��(���:���iR~#�L�d���&.����b��QU�}��)����8��DH�@�HB�^v���c*�K�̈���Sَ���� �h%͜>���e�y^��}pU� ��J ].SP�&�4�<������]&�9�����5s����|�4pR�5 b�n�|�/��%\'Pkv�t�L >�tEf�������Kj,��4�[�*�+߱{/���4Ue����-�|���/�w�̎��.A�\��uۥJ�24�M>�]�OR\�e��Ig�M�2ҷD��f�����9�񑛁q��X����[�z�O�P���I�]�~q[�|Mkw
31~��Q��[�c�������^�(���>��qTn�	�>�!+�G�'䪷�Ʃa�
�qs��䗴�]� ��\�C�����A)h��6�T^����(������)Nv�@��Q��G̯G�ܾ4"j�EW��_�H�����b�;�p�L}a���l����:'P��O{l=���O�x�Ϣ9�~ ���RZ�bCS.��΃�)��'�qz���(v�5�l�W�}����b��-�����r�q}����s�IX
Q��ۍ�C�2�O7��B��$�Y7��4O~x����<�g��*�Yzψ;�ɏ��n���=X���kF�po��Ph��h�;�J�;{�1���z��1C��[�i@���sq�-}lq�n\����[Sr�p�P��wׅq^|H�9���5*E���.��	�����*�2��uq�׺�$���P���$R�ZI	ì�˽n4����ݫ�$,}D_O)bom����m��z�H�I%�=��r�2𫾁��T����W���d*+��8#�g�|@��t��`�tA���}�p�ȫ6�u|�%/D�<�yb�пL������v��Ue���6��'e�[
���G^������3�+���R��յ�+5����2���UP#y�� ��Þ���̧�N�C�/!�u��şy�G�L�W�KC��b{j���]�<�I3��=ʒ(�'�B�J���zH�K��T_� ���'����|D�7>�p��X��@dl�0�	�ŝ�K������1�{y�&d���S��.h�P��q����xw��`�=\b�}�����ȿS��;��>g �f�˽�'��8��D[LM��m�g�^��C)/,�V4�u>Q�?��(�J�<�&�-*9w���5�4�7�㙴��"W��U;�>pن����2����A�4��,/�'�e�f��E���cR�*��߻H�]5�d=�����pL�l�����U�|�;���0�=�
7\ww3J&	�����4?�1$���b�P��¡+��ᗒpͦ��\����tE~� \Fm�P�+��O���l��|gD3��m/�Ո�k̒f���K�h�J>��BW�A����h[�&���5�^���#Nֻt�U4~B�c+aԽ	�6yƫ����v;6j��@�]�`�[-��I�m(�)��A[C0��A���OT8n��T��ׁz92c���}2�Y�'Ob�k+&�֖��b�u۪���	�ޔ���'��<qz^ۣ�̎ f��Rp��23!y�:�Έٿ��=���Z��/�3��*+�w���c�Jn����0a�*��z���\v%	V�m��@��+'�N��FA�Y��r�$7��As��(������T��3��R���L'C���Zn���=F�o����-!@@��^l�lɜ^� MgH�ikK{�vf�:�|��>2���?��q"�^{��ݭ��el�zC%���H����FM�)��U3�p��8��b��}����9v�^#��E�1/�Oa��w�	ѵV�~�2Uհ0\����e@q����DTs��:��m>!��q�M�#Jm@��6)���� �es�0zM���AͪEk�����FF���O��+cΰH-����a��gt	3L��t�~��D<�I>���Ry����H�i��H~ �0&0#�,yW�e�cH�Fܠ<T�ś�l�F���M�4{'5�CR���Ÿ�|07�P�9��{���P��R��H��%C��$���޹���Z�k�P?����ꤹ*%,>�7�ӥT�I�J��BkuO���g3|��(�1�_��j�?�c�nk����c�)=e���Q��x�b�����P=��w�-�����
�e0�瓕qS���>����	�����N��T��p�"��?���VL�T�Ҟ3uJQ���XR!���萗���G��Ddɒ8�VRM�U��M��EӺe�t���4e��oyFK$��\��'W?;�/Ӑ�.�}�Mz�Fߢ���qAФ�*pP߄bÜ[ײH�%ᠺ�.�u(~����]4||��P��yg��/�{B۟��;����l��-���t!=�!Vg�xC}N�"�ԇ�:�oH�)�h%d��Q"������YQ[��M��Sb�vVN�Y�j%��[���/�/_�І/�y�#�k��f��� gHp�3�dT!�DޟG��@�ʉ	��$�.څA��fuv'�`���.�V�z�.x.�P`�/���L��`��j�L���ņ�e!/a�ΰ�6+N>:�Գ!dFZ3z����/��Nv�r�S�]��ͦ���ѧ�&�o7�g�e��xy��3�xNsip����P�?ƒ!b��-�͊�v	=3,r��`ޗ0�ו>�&8h�\(:�̍�V G�y8J�Y)$/\� �� ��M`u��)���K'h���}�{8[�� ��+Y��}�2՞��S���'4�b̪3���Q�4.t&�Z�w>�����
UW�o�
DA�]s|�"�U#�?Qp�(b&+0~-�ٕt��8�ZN�_�Uh�u.�Z�/=RKM�7���B�17]���56u4�����2�suJ��}���0d�s��U�!�f�	`~���{{��(�pY4��yaL�s[�pn��<��K~���$�Ӓ����D�	�z��,E�Z��/'�%��,u�RO F)˜��f
,R?�Q�S��>w᱁�w4G�ǭ��^��f�h�b��<=�q'˚>�Ś��!�'̌�ۗT���"�tG�U9T`�.���o�I�~ۄU� �H,�ƞŝ&Sb�	�Mzg�3�B��F�q�j���j��3�VEXBXoP��'��%Ǟng�~8
�����Γ�$�l��෤@��"���^bwN���� ��]#�b�w�ɸ�-�j�>Gj�:(J�t��A���T3��-���+�#�,}s���gM�!D4�LU>o�� W�Fl��e��ַ����S��L��Tͨ�8����u"��g⣯�$Pgy���ܲ�*\7��CW�܅�y�M_�[<5�vk��"E�m���\l'o�K���$t�3�vlA�mp�q	E��tx8� �m�����Զm጑S��̹�W�� 9;��2Y���y���ӷ�3�NzpFb��U��Ql�;�o���یuִ
���Ðt���xʇ���01�Y���(�
��i<�a<xT���o7I�x�������8��EΘ��FjxFW�d�1�Ku|��iT�lH��΂�"��w-�N����)���Ob\ܝX�Et2�͙�rZ瓥�y@]�:&撔3�
e� ��%I�CL�I*�*s��H�a�䟌g������C-��jps�d���#~�+��S��~)��{�8Ng�k��pj�"�����U���f��I�:��Fɣ�ΠH��inoC
lǲMN%�*�6��
�_+N)8Oezw%'艻U%�t���x�n�z���ytH�L�O���-�?/��+n��;T���]��yV��"��)����?1"�����Ʋ�kQ�P�x�T§(���ۚ�_���:��Vz����B6����5��ѷ�r�^�,�K.�8��#��J�?��65�>p#W�6��$�Zk��BzoD�#�n�w �/8Q'.�r5'�h'v����,e,�\����V�W��y:
��Q��3͢�Ԋf�LR�	<g�n�H�j���@�n��^��0� &ӟH��[}���?z{��� ����]�T��6�l�IF�p�p���!�ȵŋ�[�[.+nY�h���8m��^+;�Z^	 (ї*܂>j��������{�%��
���,T��x�}��y�{i@_���Z;�E4���~�/4Y)��M6���m<Y�ѝD_���Z�0��TT�o�I���zd�_�1\����3�/����7z�v�"�H���r3T+~&Zi���
Fם�o�=�S��5x�e�������엍fI�g�$��ivQ(_ߘ�b�ߘ�
f=ܳ�r�Z��v^X?�0��7��8��IE�6����H���)�%����8��R�>��H�:В$�P���
�ikEN��'�.�l��_�>a	d�&փ��Y��k�۷s|��1(���=G�"o���]���.$|�7�|%��A�+��3�h�(�	�3.a��EJ�~>�� ��gj���h��h#�x\�����P������kF��"jk/w�p�T�[
$���_���Dn�g#�"��!�l�JP|'�-ˋ��ad���`��!9���`�>��j6{� PɪJ�U8�-�A�B���U�l��`̢qG�+�n�a��]F�j���[�^�'}�g���
񁝫�����Le�p��������Q��+�8v��B���� ˳���I�$?��	Z����JcF�E�ҝ�͟<��e���n
h����K1�l�}yL�owߒ�az\�S��B���U9�T�RV���4͕����/��u��Z���c��y���A��
�*��g����b�ǟJ"DKe�#�=e� �{�Q�	��Lo�JvNo�bs�,��>d��[�zd��ax!zs�f#�|�	�m#5F��h� �,If{���2C�t����"gx{��eu|�����qJ̬J��[�FS�^� ]��]簟ļ�+��|Yٻ,��U�N��Y�;�뽲7�E�Գeq-�����ԑ�0�0��I2~T��cL���q��ԅ|��J/s�t"���۳@�3�6����jӳ_`��n!�iV9d'u�Ю��Qv�P�:�؈�k��ïR|A�U�}A~��4#�.�\�9��8H�~M��
�muH���Au&�P�
�!����bWk?=��:����l��q|>6A�D�y:�D���&�j�aZe�ɿ�|��e;:� Tt #.	��	y��§F��ҏ&�9�_�X���+Q�ز'A�N�����U9�k8��3���'�u�_�Xa�"8�#q�z=3���<w�uVը�;7<y�GΘ�p#1�	�;��L�Q����=��^�T�t�)�	+'6�Q;���Cj�Cu1�d6����&b.+������f�^�%-�\y����7
�`�� ]�,rʡ�������$�n_ؼ�iYZ��g�: ��d��w�-���U�mVuC�D�Ax��к��?�@�/3�%eB$$v�A�ռ-X�6�f8��e��F��R�<��Tzy��pJ�8j@+��G��JX'K�ň�%���y��m·��i�3����a�kV�җ%h���: d��<���4�s,u/��u�N p�S�8�.7���G@�\���uwS���F�P�O6I�ī׬��*)�ލ�$׺ѫ��%У����A�"�VGEC�T���<��#+�K�$![�.f2g4ft�
�Ϡs�����%����w��㖋�i&�Z�`,�;<�*0R��u��d�m��%����2�b�_�˸F�'}���Z<�#j��NJ�Yo�K돴���Lr��1#ʆ�<8II���͇�X2�K8K��.+p-2�^T�hQTp����O�0}�~x^��|&~�����,�o�
Y�P���!�;8謾=I	���Y2+-�|��Z
�Ǔ#��$�&c���������D@c�Q��z7T��gt�Qk!0�8�%2L�F��I��T.���Ԋ�}��"�#O�E�Q�P4n���eUO)�[5��#�yk!�M���%gP�����|�`x��w#0"��pJS����d���`�R���ԓ��l���A=��j���|���~�Q
��P�!O�.h��ʲ@h`Y��?'hͨx���EH>��w&>;�K�iti��1��)xw�gL���G��Y�E����oC�!�{�ՖkĠ/.o�����EF�ONؙ���� �0jK�vqd|ǥ�六R��j�A�i�v*�E�QK�N8%�9�N�,{����2؜�������S�8�l���s ]��P5pnK��VSS���Q�}3�L4@.fM�u(��4|���M���[��FEI�CO�*�-p(��/�E+��b ��%��q���-�үj�,P�0��QDf��V�m&��(�8��F9�iϣ^�����3��1�q}�����?m%Nvr �E���1�|5���-�!��|�)ZUN�T�ŐM��%֗pn%�=���ГO�XT7����C�)^.͜)~�\�V��pL4=w��~�)*��c��)%0��t�XP��I.Ojw@LёU&�rz�hW���K�E��Ǽ)]�jb�դ�Q���KZ%�k�g����歽���@�*�6�èl��>�^#
YX�����ƀ�&pb���=(���3����l,bŲ �֙9�|��J��N�nl��06�P����[r��y��;�/D���7!��BY���Y��Rv*��f� e|�Nc�4�h%,�^�&9��v3~#h�6��b�f<�[�����kM>
-�7D�ń#���7�u*SҸwI���T�%������)��_��l���ϋ���\��ٙ�����lwa�JY���u"��8'�`���+x��v1.Rʾ�6I�K���s0��e�����������C���HZ�:�![S�Z�/��&I�_/���$�<?PX�׃c��lCЏ�nۤXk�<;�cV�_�H�$��V -�����/r`�����}���W�!���G�A� �Ío�/��@��4qx����Y��V�;n]+�Í��i��\q9�kSW�}�&'Z���-��^�N�kX���?.XhrcQ �h�4&/��)sU�܏@��w�CS�Z�)���U֎����SW�����|��K��`�� ��Y�_���@�_Љ{�)��bJ"ܠ��]���^CP��R��53}f����G�M[�o��L��<m񳂪������%I��v7��|vzj�?}�m�2���g=6��r?�ᠭ�p��Q�Q٬�y���N���e
5#C�ʵ�X��\�G;)��%{,>��K[��+&W��#�1eL\�	w������ݾ#��gi&r,��>mz鞪2��g^�`v�z�� ���>�Od�n�.���x;2v�P�9�]�%")���2��/G���Ȁ|A�?�%ņ'���b��^h�xE�'>F%�3&��s����̏�z��c�>���fi�d�>�+z�	u�J�O����`/���]��G���ZL���m�_���1��׺>R�t��߅�SA4�Q6���FmĿGo�t|c�ןC��c�O� ���H����s��B<�1�,7|�"�����z^u:���ՒW�	���<)v��d�k\o��jƘX�VN����6а��}�=VLm�p�cb�Ǚ1�2I;����ko��:\N�O�t�j��.�W�5�J�s�1���G�����<^*�j%S�s=�e��w?gҘ��ǅ�|`6�8JL��\8���@
�6&��^У�'x>�fW�y�|䦋���W�A��;��|3�*	�k�S���7�>�{Lb�AƄ��bQt����&'w����[��
6Fv�p�JW�Z�f�:��a�Ov��W�T�vrA~¡�i$Y���K}����:j�^tu{�U�W��/��?Fs\�/9�^1I��C�&��U�J
1���<R�Ov����5JĒ�S!��L�!�'I���Y+X/I�kwlPs�������B�� ���E*��E(
,Mo:�񱇯S��!�Lp�I�y�$�<�Uw
V𵇪��{����ZR6&O�d|�_�(2BK�1%b~1��������_네/i�k	��"
2��L�� ����/,�@�^���o	���(�*�'��b���o��	���1~ ;��/���5�[�����i���r��P���1�m��?7�)����fQc�yV��=��[_�&`>W��S�����ڂ}�t\�i(X�`#�3�"H1:1��p��|3�]��/S�u�u?(z���CƋN��;�H��b+�P?Kj��xr�G��H��#�w��$i_�q}��Dz������7����Ie���X��]8�G(�৚�w�F5����@Ӷ)�sB@�"�'��_�q�����f�����i�qSk��A,�p�/4�/Dz���/�-N�}���e�nn�>t�,���Ou�l�]� RݖLs�TUXtX���ϓ���b�ݣ��r���P�:��l���١����SN�� r�*�i��sp���>�f����*�3B�6�'���u}m�p�zh����wo^K%�^�nY�||��GS%���� ����4+��"������^�Կ	�?�=��˔(��b"Mk\��^�>��� G�2��B� ��_2�Z�L����E`>j���f|C�Q��=M.#_�;ZҞ1��}���8�ȭ%��K=����Ǥ ֟#"N�ф�˨f��d�Ź�#z�L[�m��m�m$�=W���-غ� v��l4\p�������~�i�R�_���LTH��E��8�0��oh��_+m�AX�<��e�rt��Un�3��(Q���5�[��w��&��JF�Ypz���8��/t���;W���=l����d����M��	\@�º��8}�YS���E����`X�QK��d�!���)�Ha R5�ڗHW`�d�������?d*���Xξ���\v2��S$�Q߾�/f1]�E�۾�.���7Ś��t�Bg�Kd&CۘHa���V;w�z���Y�c�?�/��3�A
]�8s#�4�߶�̳5���"�~�l`%�Q�4Re3���لf���>d\��+�kc)j�	Dc�b�FJ�!�C���.��69��ܫ�}���~����[9D������sv��u����\Z���X��[�1.��sè��}n9ϵ�9��D���ѧ�y��v��!��>�J�<A��φ��NR!d�r����#�ʑ���}�6�
M,t�E�n�,�nl4����Z�t*?�~
��=�3]`|P1�&� ����������g4�n�O�n��SS�Q�B�.ʰ�X�VH��L7#6	��y�z��E�I��Ձ5<=?�#��C��^�E��@6�ǽy�X�K�a���BK��Ţ;�{�t,�@���,s��rW��͙+�� \Rj$���6�W�#`J�l�U,��g�!�i}�B����������fHc&"�N3J���ы�-d���n7b��f@E]�̧���/·\�kf�PVtCz�>��&ț4��ɐA�v��b�oeQ�����XL��|�-� ���(dB��8��d��k�'��J8CV�u�Bf�޵���_��l_�NS_�h��h�G�5[��5<�z�4r"�N��h5o�X�^�����ޜ)oDeKq}��+J�&�, �!��\�a�O�]�
M#����FOô��Mb���4�|�C��hA|�s���& ���m����޿H�
Im�~Y��
���xB�P,�ruCE�oZ2�:-�xG����):R��NxǶ1d�>�:�L���.q6;9ν��2*O��.���L�D�l3wz7������)�
g��e��|�
Ǐx�xg�м��kل3���I��@l��Y;�
-D'a}d�h�?<bqn��}#����v�^������\�?��?ˈzȬ�Zg7���g4�J�o�(�qo\A�>�r�+ǱÏ��en- �+�P\H����U62!�j��a�U!�����U[�)��#��4z�Z�_� ��&�w����mF6}	�\	�-�^c��WX��8��)�������@#/��*$,�l��7�u�����R��)eOfQx�D�`�E�d�,�kz�c�n#O�:�&"2��*,��Y�9�~�6oL?=H"#��.4�ʽ��4�z��ڛC�X�0;A�e������=�<N���!>��G�mnYt�C��p�L� ��*����m�aϢ�P��z��e�SEy�hY�QH�U��ܫt]j��ͳ:�|P�ఓ���w��O�q�]��/�R���_(�Y�}��&��>����t���B eC�8b�5�a%��r,	�1� /@п�E�G+� �n!�� ��F�F��N��"=gq�>�M������v��dj�Y���J�M�<�ڿfdv��S��ƈk�O�%�B������M�,bNIH������J�5A�l����Qjz��m���Ә�s���*l��7�h��|�04� m?P=�X����R��v'��\M1h�>�kk�}t�_mjSP�������^�z�и�AQ�V�b�ɰ�6W�QD �Z|�b6Ρ��>�����P闔���O���:�V�
�g {��Q�{�}���M(��~؂��2���NK��T!>�.�"�W�%ȏ˫��^���~��+�A�y^b�+���whV����������U^���*����^#��ɗ��N0���}������Z;�D�E�-�%���m���8^w�I�S�%��F87Rn0�&[��<?�f���9#��Т9�e�s2c�T��e!dR3� =�@�p�"�V?�hc&aJx�'R!6ѧ8e:����

0K�R��V��P���L��<$�nda�&U�6�Y�p�@������"Esl�G�*��m=� �NLǃ���m,�F��3<�>���Գ C���=:�Vup������1�6���?�L��[+n�4@��8�����gVz�c��ҏć����k��PWae���{��hR6K��M��V�\V��%��y1�bP$��g*�p�|㺌؁�S]�� ;U��`V���X�6s�ȋ;~Q�'��9~-�z� ��T1���2�Рŏ'�- =�$(=��O�\V�ȇ�C�̽u&G���Q��a���Y��9��K;����3�xz��уr��,��3��O�2�Ju���A��X�+�@�����$��í�\��@�e����T~iK)��|):�c��x��T��L?�AZG���jb�S|�X�τNc��	��R�(���� *QL)��e0|�AP�쮖;��E�.�O�j�_����FQ�?�H��K��q�qJ��;"��x�pY�dK��vJoD�#��8	~�`��]`�b�N��B lZID�a������"J�w�{g��]Ŋ�B}��Mh�h�37�a�99��\L�{G�a�͆3{2��`j�0
�D{���>b�&����]�Y^Y�iU�sCz����e�Ϛ�*��u6�3�≣ԭ��u��(�_��WG��<dܳ?$�7���D�n��J8�&��ƫWT�I�=�������MG9�	�B��υ'5�;'��3�VW�_ΠU��G�S?n� �T���6�Y��?��V1������",ܣfA��n.T�� ����N�m�ZV�*U��k�"+�"z+������g�.�2��M���u:�G��	zw ��a�`�k-��Y�L9ʾु�l��|���Q��Ld��'�+�٣>��o�� ΐŁyM��4:%KsP����tʭ��T7{�<QD��V~"�A���?��e�� S���1܍��n7_3T����F�u󂴏�"9�KsZq���lwZڈd��G����iyeZ�؆s���r��;1 �P��`!������ܭ"�3	E��!���������i�%b)�)��U
j���M(`u���A��U_��c�F�
?R^	u�7?x�н�<�~���h|�G"?nS!�ƙ*��E�o2�H�����NF�pax�G�hM4�S�9)�]���1�����jʖ���Sk����х��ע7�b}�q��Ϥ%Otg�q�4sEy�V{g��c�&����\KH�{"��A������.Z��T��N��
X��I�d�l�{l�䙸*,=�b��KKe�q��;�ڔ�T�D�1:���LU�
ALH�WR�D��R�PK�G�cKF6�Q�=Xl�³�e��-~a��S�.��
�6����g�C5�F� !�͗�R�4��=�+.����!j�� =�Ts�@���� 1�E7B|D4�8�&��{E�=n�2� J�CNH����,����">���(X<0"��5>�϶��۠��󅁭3 ��2B&�{��'YmVȕ��u1��~�W�_�?$��E��}���Qe�.,[SL��C-XST� ������������Js�AeI��;��	��0��{".*���
$MQ��I{	�0&��)Ya���FY�����R��x	H��ߔ:��3@v`�Q�he{�*�<�e��	
�n#&�l��X�R��G�>����lױ���p�9B��1 A�̥nS��⽨ߩ�j�9�2��_��X�	E���xc�����"�0��g�Zq�`�j⧗��T��yak�/-�f����^�;-�������@3�N>uC�{��8]�32� �#� ��c._��G�C�X=�s�F���&����J��%��7���{̡c�3�R���)��]��{�*���PLy\���AN!�O�� Q_L\�U��>A˺"t��ݘ��%?�$ugfjz�W�� %y�ߌ�me�	��\aYQ�[��N�"�6@f<��3A��eP���*���(�vN���9R��(���d�Ց��D��aC�/M��As�g�r�R �Lh��#I+����>4�x�-�����\�ژ�QN�����<�7���:�^�}��xn�e���0G�oj��heܴL+*4��FJ�'a��4+n���Y`���>��Eb�͚�ʮE8�aG�Ōʻ��s����D�z���h�FӨ�d'�����+l�X�M�b�t�eC���bqm��.~�e�F���J
!`�n���0�@�Ih1�=��g~L:'�����z�T�l� hsDNС��^eN�����S�����Ũ�g�1[*�e4�4ˮ��!����B�zu.
L����8! ���(@q-���k3%ً�K�X﯀�������6��*n>Y�%��ހB��������xت�Ƴ<C�Ck�U��7�h��`p�J��Dt�'���]A��U���ȴ5�=�<�d�-E�E��(LC����l|,j�5��>�G� �N���j<��V����4���h� ���Jm�,Xde^en�1�?��a�=�����#�i��K��#�;fD��������r��pW�,	:U�/� ��aG��#5a,;������F�gᖯ"2�d�@��������"S�g��i!�� �ݣ�S ��|�m���4{���x�c������T3��6��t����=�Ǭ� s!�?5� �}�}�W�Ì������S���1��4R;n�� ��o��@��>��h� �ş�����<����i���m�4~ķ�h�����?8��wLN9sqL�haa��aXu�ڽ�B�a����u�p�{���3���eA�������3DI[�
* ��xy���f+]D��Jl��xD  �X��������]}R�}}Ic��ʥ*�J��[���q����Y�`cN����KK*�����2�GGO7� Wxc|�!�ǝ%7a�*����Z�M��ح�۔��ׅ����]���;o>sk� M��� *;���w�a��=��p����G�Ox��͊^࿿B�}o�7?�v��@L�Zׄ��$�Ifc����\�P�!����7�
z�}�T��˸�e� /'�)�u��u�B���ly>���3�鳯�p]����� �xi����<K�O?�O��D��<��r�"[�i<�Kr�`�/���WS�O,�+k��Z��p�SL�30��"*�$�ʫP3*�؁�Y� O8�p���Y�03{H�K�@�,}_�~"1�̓9�;�6�n�  ��?�K�#�G���dˑ$�?Lo�m<���ِ��������?���o/���} �/��ǒ:gj��8}S�/݋��WI�痑��J� }C�� ��'��P��4��3�I���:��� S��qA�ȵ|�۬fOP��f>6�2"J�5��)��L� ���	%v�z,O1�>Y!���2h�""���r�JH�?WqB�����m��a�s
t���e�.��O� &~�MuR���ax�8	]d�c^Щ�g��Fj�-ш���mC(G��1���:i�[�W��
`�d�����{��R�q���8DJc�) ���3h�.�fd�$&/��s����Ж�4O j_�b�92v�f �̅H���<C`#g'�l�VwS�h�!�eeL.hQ%��j� 7]�v�NI��@>!�\_D�O� �S�Qچ$_h���F���N���>��=���r�3�;DJ��J��u��ߒ�C��0FΩV%�g�
�]@v͜�@����c��n�n�F��
v��M�(���:�Z,�b	4��G;���z��D̪�&�J:Zd]ʇ=�p��������چU�R,��.e0\.T�d*v>��%����]2�S��p�j���B�G��!��[����o���Q���".�щjWBp!8���K���C���,�� 2���O���_x�|�5Sf�������)�=�K��@����³�[:?�%���*$}�#�	�l`�l.�>s��`��D��h@��4�k�2���Jb�F�Dpd1.������ �m1�T��S6��hy�*n 5yz#�g��'����O�L_�'�#9��/kI�nٻ� G�G�Q(�J>C�y\L��A�fQ(��(�J% �r�{&cJ�
0�l|�$j�,��EH�:"�	͎T�0���_�(i���~�����b�3iW�j=p��/�� ���c�X����h'1����j���p42��|�	�7�$�1�EMJ\Ѭ��� U�/�~a�fӆ,L0�� *Y�;N�޷�f*]&�5����������Ǜ�bc��S���m���ZF/�:��_��eؔ���:����B�2�]�M	�����?��i���X_V�+W�7&��f[x#�� (H}b\�����~���ϔ�A���q��b�0/:�Qa����KB3ߝ�>�m��v����N�L(�(XҦH7���j� Z�}�X5�7���k�'%���8�}�����֡���K�[���,n3/�6F�'��n�gm��?�>�/�e.���l�h��[�X�cFn����qo9>�>��1{���^�m����4տ�r�����V�����M�`���ҡ��s��>&��(�0N�M8V����{C���D	��mL� N�x�N%��Ϙ��Yoi[�F�=�O����W3c����S���~Y
 oK���F-0;��/~a�R�gq=�ц�ыJ��L��Z�T0]p�(�M�%��F�O�Z���������TS�_o�,� ��L	���?��A)��^n}Gv*��B5���L) ��N�s�o^�\#f��<F� ;��&�c��u��* ��.m��̻���� 2ǜ�Dֽ���\!�C�9�P&���O���4�7��� \oC!�`bB�t����K=�%{tQ��?�MO{i�f��� r��i��X�.-��m�8?�.��SP�?P& �n<��id��:���O��&dr�0�"2�/�� L�c9� g���?��Iu�P����#�7�/�I�l틭�P�N%+�k�� 
��W9��}�3����t2�\o����	S-b%�	�x�t��1��E��9a��{�)5����Op�n�~�
~z�}��e9h�@W��U[>�πB\]�����uk����!3m(~���
��6�9}��
R�Gi�~k3ڍ�~�I�9S��W�%�([�7�
X ��l������¢��
މζ24M5I�1|l5*Z��>��3�� 2k�~g�L��?��42����8jl� ��\$�>���D�O(4J'���	I.�+���x���K	��;'����� U�$���@
q}c������ �_��2��|��c�\��@�?^������~��1o�
����4�Xx8e(3V.��I(b�L�T��L ��U}�ёqӿ�A���f��1�s �A��M���~��Σ1�*�[�+�,�c�X'��� ��%HŴl!m��� ��� [,�O�}�[8��EZja4ex��[�� ����+(;#��� �N�r���l�e{?�y������YyG'� �)���%����+�ph6J��+A�W����ޔ��@���~yT�z�n�+��b�-6Y�C7"���L����/�h�Ϛ�+�Kѱ)~HW�@x#���߄��v q�q�/]�B$hT�l/�!��)��Ox��p�I�#�(Op-�qC�����C�B�/����TY���Y�]��_#�ŏ=�#�3�k��~譻h�S2y�6���'I�h�Ѓ�0��h��n���.�@���q�J�x�^�ݡ�
(���]������n���N�QA�W�D�a�W��-
h�L��$����2��N#$��S��lp����\����?��h��P��RS�bb�[�d���8PY�CbdH�	���✳��"`;�� ���#�����I�Dt"4q=��ڲ�F��ȭ;�oOe��o��c�� V�����
���sI�eG���x���GJ�|�u(8ο�FA�?��r� k�����X-Fa�X?��O/��a>� 4�=���Љ�w@��Q`�1���� �s�3�W`�܌"��	�W�P����/�_�L����!4�� �h��Pc�N�jb�_���6�lK�Rn*6}cl?��M��]54c1���ME����eĵ6� ���W�T� ���z��A�Y؍F,��D`Q�t�\���5�	�4��O�N�xp�b�?fŮ6�K�J�����	E�~h�@�i����Bgc@]Gm��;.�;�� T��տz�O���P�/P�B]�hJ�
�L!��!�Fwg;���c�v����čWM���pbs����8�<[c�VH�rH�?R����t���cHW�N�aǪ�/�� �Y��}C
���u+,g����������z�jPC@�^�2�e-a��G��}������d���-x&T���7������?[&���{$5n~��{�P���ʝ��O@�0 ��x���"�k��v��v�^�<���`K*d�h�z y*��֫��b�����5.� ��2��b��e 6w�:���֪��%	Y�e��j��P ��&4{5�I~��Z�_� �n"�� �k���HW��o&��H�!�)��}ʰ��>LP�A;v�l��ٕх���W��V_��HEv�eVfc����VN�>\N�nx��X�D/��z>"� 6�_ ��D��G�5��~�%��~��������';��ҝ	/"E�-�+ԏ�Sx����X���v3	��'R7b(� �#�=[����`����+�0��; ~.�U������eO/\� 4�����K`�ߞH�j肢8>kD]ZNty� �1������U���El��\n���p6�`*�ݼc��h(�O��.��YSu��j�� �'���*EE��z��j�����:���\����c٠��G�W��D�z, 1����Ŕ)����c/+O�!�"	N�.�<��~ ��NH Q������/��x���BYѸ��[$͝�/��K���F������?���ܱ�ɉ�=��dV�i��P��{�_y�}���#1��؎U�G�x[$%��&U�/�/�O��g�c�V�e�WX�h�w�P�޿��3rfJ=���"��!6�+1�p��T��� 0�b@�X5�Q=S�!D���YZ�0�yh��CG�P-h��I���'��-���FXu���+b����$�`�V�T�bB���p�r<>
P ��%���%�l�2��$� <͞7L�d�K�p2Y���#���C���j����DD�>4�̫�%X�l����0_�5�����n������g*O����ss�g�9/4IEj��Rl�`= AR	�T0u��0h#�P�e����p�i�Zu����N�ݟG�&���>������� 8�/�~_��͟��cs���m�y��z��0vkiE-�HhE��CpV�29褐d}�� 1���=2�)~mܛL���8��mi M����#�Q3���x�?SI������5�f�x����a���q�UYB,���0�w��	Ra�ΘՎ�� �Q��zO@xW���]1n//�^n�6�3���������� >3Jz��Ot�F�ۗA9�=��j]�� ok����-�u<q�r��eM�T�ځ���0g��A��U�Ka,�Xlsq��AX"�-�,�X���4���T�[���7F��DB ��}��0B��]�K�#�� Q��ˢfyA]��%(�؄ Uļ�[�h�^�%�:�1A����.����^�W�d��l7��9�F��COࡈٗ��Wݠ�cK���-g�	&\q/DO鬈�Z���D�0���;�V�,�Y?a���Ŀ�t����*�yC�Mw���o0/�[���&m�Śߪu���V� �ο>L�"'���N��>�-��0	��X��&�@��<��_6*�O��,�Ѳ6�g�P%c/��mPQ���wG��]@�}��� ��CLF��'�[١��|`����y�?��"J 0	B�V�p�d!v�!���J��j�!�ʐSV����`��σ�Ӄ����eS1����{^��� ��«�W+���R�*�^�>U�����P<SQ�<FaP}���>K�8j^�`��&/ۈ��$�&)���G���˼����ڿ)��p_�����~�/ ����_C/���ۄd��T:ihe������b���@���=5���/�,��뎹�"����2Cl�"}�T	��@��<���NEB��(�=�=\ǡ�ٍN<|�kE�x�uC?ˀ�ao/�A}5�4Y��yº���P[�Ǳ��%	�0g1KF� � �5Z'&�:F��1M���h�*pL�Ez��I4<z���@�r;[���s��9c�o�M�E�P��4� �#��+YQ�@l\%s+��;�Ϸ���q�xTmB�I�.Ko#oЍ�5�(~*&���~Q���g�1-~l*�	�{��!��~C/O��4�ڛ���Jo�+�y����CB���5|��=vK��gKe���aQ�l�u����;�^y�h �Ͻ�ɀ������0�b�6�
�k8m�u��*4�O�!v�tf+�\ZM:���`Ò�;����o_�vը��H*���_툗�Я���+��wZ;;vK}���f >�o9C�G���.\$.��.�\_�kN��Q��4���9ڍf���u]��O�0W�'!*�&���� ���d��� P���"X�׃�_K� Pԧ&����_L�[�� �� p��ڻK����~4Y��O�o���1-�B(\f�F��*H;1���g����[Y�g�PP�1��zQ|�ב�O����-|D�Z�P�oũ��~�;fA;���2�A
� �u̐��B�}� �]�^�d4٭��U<~�ѐQ�W3Ipy�ꬪ��u��&FY� �z���J~q��|>FQ�TIB� �â|��"�,�	c� �1�����!�O�収	��P
���������5��.�ZiKI �|ʮm��{��
��C��G��W�S6�R��t����hvK���F��Q������]�>�Ŗ����_�Ķ�m��+��X5SݰXv�WTaz�v��_�(p��~�� 
 >:G��>L��,�Ր����#����}�����_�2:7���  GG�Y�
"��~�d�P�k��Y]ȩ�uC8��� ��Z)z�LT���+}bb�S
�qK0�>%���}`(�R�^;!@���������l<�����`�e0���:#���,��Vf[�E�{\��K�d�=$�#��︼��A�ql$��o'�}���ɔ��A�I��T{�|�rOf����
��U� r%h�.�ȗ�(Z�P[�E�2�N���oߢ:_���
�Y,�w<���|�#�w#�����*e:� �d~��R�s��{�� �S5��|��ssp�b��P�f�10[��w���`�g���&��*��O+�s�����'A�/*�����E��>D吥1�bb������[Ao�. ����?�P�bl��{8�3#�0Y�<umǼ�Ő��#�t�D��£7�0�	4��
�[A�O��R�r�����, �ݮ`p0�&x�	�:���nާ3.d"a7�t�/��1Hmv�����#P���ߊ��#$�[^\��5f�3�p�"�q��(�Ř�X��9�xVЅ;�~�aD:^&����؁@r�J�/DET� ���S�=E�a�-si��a�Շ��h� �s�������˔� ��/�~?��0s�7�;?l����(�c��ŀg��i�ARִg1/��K�X=Y�)�bFl��v�3�wAq#��C�i(��w��t��9@�<�F��3�eN�:��~*tC�+�<}	ORV�W��xpDX{%v��J&9��#ph<~v^6T*��Y��D�Q�Q(�J%�V����e*r$�CDy7Js�������փƕbeGĽ}2M�� h�.w�eH�z��9������%?Cg8�|�<����n�FX@~�\�*#��>���aG��Hi��D�f�b��c����,oza�w��m� %5��_�XN�h�W	�x��{B�q�Uy������_�~-��)0�M���2�96�f����o�۝T�"� ���I�}��-�Q��<��� �a��'��m?(h��:0%�VG����V�RU��(������}�@��:�Tp��~�W� f?2:�1/o�0��m����h}cO<��C���4�tT����������M�M���{���3d�������bƇ�G�Y��-���  P~�ߨB�vl\JTi[���,ݐܧ�K:ћ ���b�I��L]��o���<pB2>��~�]e����	0b�}���'�ۋ���п�����K`x�<���͵R�GYR}c�֬&[J�v`!��l��MN���'�<�'��}>��>SBI�> 9����R-�l���2$�>�0s�|���t<%�U<���NnK=�q~�A�����퀮Ur�^���1/�&ue�mre��Xb�@8�a�~S�f� #�y�z���L������h"��ae�x��:?��K��l{ɺ�� ~9�[۴>#�M����P7� 
>o�.\�4��j��UN�����1H��j �����c2�!"�'=KR���})��@��0��_$��7�V��D���� ���}B����%�OS����q��ɰ]r����o��t��b�}���e,�7��d:���_W�K��W'� ��&wϫ|s~�@Z�L� ��!�Uiq���ޙ���$��{� ؋��j���O `%?V�O��� ����?�a� S�/����|݄�t�,),}������?�D���=�C`��3� v�O�83B�γ.�D7��p{;�;Xw��c6��/���S� ����Ȟ��MaR^%J�ѽe2���<�<dW�x=�����t�	`���g�_�fn��J �	���/R"��b_��3%J���i�Ã>�y�v�=8�jg����M@t�܄௸@�>����D�LM${e�����"�)��[���)@D�j�b�Kw7��`cR�����>�@�����E}����
�<ؒ�
E��r�4b	�<�i��D9	^��Z�+���W��f�/(�b_1��\_����*���sN�@`J}>���e9�� V#CvǇT[hO��3C���dyÖ-VK��ԫqї���_o�X�#o����g����]C���dB8�P�r{2n	����@��{�a�ELL �d��a�h@����3<�(�z>�,4�$�o�4G�2 �`�(Mm.)�`�p�p-�Co�l�\,�k���*���
(p�U�� ���z�u�a0b�����JACY���.	M�"��,	�y�`��"JT��Y��%(�B�(*�hƂ�:�H�ߔ��b �����1�DG�S*��G�	����W؃�Q� :�0�D7%�5Z.Ș*1c(=ύw������ʞO�NyܽL��;�R�[��,og2�ksN��<��u~�b�����k��ϬG($2��� w*�]�/���ѶD}��PM�;��
b�TX 	�c���T�ޠlkB2�jX����y�˾�U]J�7b�`F��ޥu�r����Wpe&�x���"=�1�.�v�����#LM̫>��7�n6nكIL���
\ND�
�����Ԋ&�Ce'!��sĉ�����6!�`%�g�G�U�&cM|��I@�-���l��b���R�5����U���K�vʃan䉆�(S ��`��p����\���y1}�=�ѕ)�q���yp=9f����+�!Lx(��ƚj�s�m����#H)���ڱ	�a����w�r�m�����h�O*�3fҵu���l,i�����<�Tbg>�g�xE��+}�T���#��d�W�<�7��p����s1��5���|DF�2� ����#uu� [2��Q�1a��E�r�k�F���|+�(��R�p1-�)�a�Z�9g�2�ť|E�����D@qd�w�� �K0��E��*�7)VFs���^oÇҦn�;̀�z� ���-cS2Tc>���r]��/,M�PTc`��������C��`�`��J�2]��jJZ3�
J)v����.63*3(ӯ�� 
�K��
b��|�<qtE��RS�cq���1���z�EZII\	j�du����j�u���2��!�lbY�'i<�EY���rFl�9M�b%D�,��.�}%�͈��3j���S�k'�&+�4Xe��XoQ��\�-2+��虣m� �QW�EF`�1x�U�YN��P8cG��d���@"wMK!8�A�N����	��r�{��&�9:��L0[�E�M��̏���W�BE�,y�p�y,V5���#�i}���f�N�h�ᤄ�G�L���������[d4,���J¦*�������-��[u���{��R̰Р���2�w���~euԻ *�� !p\���_򊠼�wW1 �D�c.r�tQ�wR�	s�-���(��,<�Zx��\̎`!B����e����,#�#�|]�E0�Ex��=e��3�Ⱥ����⥭�usc�>�_��V�2ӕ�8�Aڔ��=��`�x�9��s+w�B�>�n�i�d�wFH|�pKN# �Q0�Z�Yn��r������.ś20�����[�1A��:$QM��l�~\����(��]�%߻�l=�b�\�V&�|��~tU�� (�?�iE�)�P��X�6R܅o��Ǭ9�J�Ƣ�f%`�T.����� D��DW�S$��l����wd�įR�H)�X�^�/3�l0J���W�&*~��]��yu�D4�:���`x������c1�ݗ4�R J+0j�ȅʖ\+(�����S?x�}/+�\�8�x94҅߼��}ARq-*�㨡����nSʤä�=�Eo�Dsf�8<����4ƿ`z&�]3U�D*�t*rn #�y���R��{4K�e[�����TXy���pŜ|3���*�Bf䰡ѭM��ҍH��`,Cc2ݼ�*7��`��	��LpW���,J��0aqr���R��H��R�;��Q���,#��-��+��C�/�U�'V���ZhQ�����D���\>�P?kbR�7u��ZK�7RR�@#��d��_s*���e�Oj��H,�[̾d9��K;��K�ɉ�Z=�3ws1J�c�e������S���h�����[�\�ۃ?�s�,�XU��7L�f �`wQ([/�[b���K�W��<�ݔyf7C��n��~Zt�l�[9�]�U�;�
��W*�D,N�q����4�)�Q7*�����;����5�V�QQ2�7+KgP���U��b5�&}_C���od�)�}�jn��%�b���Z���M�*/�1��PVʶ�݊%�q�$�X(��=���S�0�3�/��A*ڍi�<=�in��W1�,�	�<���δg(�� E�<��H#1B8���0���q!Gj��A�o���a��FBj�X�4xT4�p�u�<0VQ
�i!�>ȍ%�����q�6D��Ԧ:��l?̽N��͇��[P��z�mZH@��*�L?Z*`�����ol�j��׻�U=�f��B�r:�,�>�������l���:�>D���i?�5
��̰]*�h6K�qxz���~<�w_�r��u-�V��
<��K(�=M[FȖ�pd(A��	n�ِ9x�uTjh��՘�߈-�t�sB�D@"���m.��J9� �;7/��`�M���"��x���r�-v���&ڂ�+]��uC<(�@;����R!H��,>G ������Y8��&����?AU����5{	~W���s������"t�g����}�� �O��%����$�.Zk@���փ�B�\�޺�u�]��6	v�Eε+Yz�.��?mt������{`ҩ�n�мi�ʃ��T� T5���R����>����F,]���0Ď�Eԭ�a|��v5�$�XPm�48�U�?p�H΅�,H���ǡh�N&SH��,�L�	������b�K2�2�n}ODW�����΢������f"Ͽ� ?��P��x�'�}/��iP����k�!�t`A�U�g�����hY7�_Z�Α�1�������B��L�I�n�w-[�d�mtM���8�J��	�C�)�l�A� �"A� }�1�;�eG�'�q:!��/H/�Py}�F�-9�s7G�o�����Atz& ��R���.i��@�f{��ס�����,�}�x^� l$�� �LBh�䯡�n`�<#3�n󓁸h0Z�������F9�*�R׾5>�����g����\��ϣ��"�^f,&G��
= @9���Vٷ����\��%s���}������jP�lĹ���C��E��p�Vot���Z���0�P+娭���Dx1,�g�����\�Y���G����F���Ԗ�S�}ϵ�����[%.tz?�/J�.�;Έ�#Ш�O���eK��oޥ� \�T���>����R��� K\�G����>�0�x��j�=#܊���5yaO:����7�).B���᱖i��,"��b��{��L*�;�_������,�u����ƽ�	�{�~X�X�=���VX$����<�JDe0�3?���t�=2���aaZA[�'����/�y^N&C�z +�	w,��K-��	vA�CS�����{�_�1M���t�\.�=n����c�~g��WL�����J�b]zV�NR�{$vއ��/�:�s� m �?����*)����߿��XGЮH�  �z��1�b
P�&.����@'�6�S5����L�M�m� E���,,E��?ݷ�5hp �t�Tl��>������d!R!�}��=߱Q5�!�cP��A<�؊o���*�� &����lw��~�*����L�[}�Oh�@X������Ju�(�J���1dy���R2��(fTa����"7���L(E~�f��2h���j%�}��Ǵ0�!j��ף���|T���u@�]��t��j�..Ⱦ��������Zb�� z1�r ^b
��o�=�!��V�s�=>�T'DmT��~f!���w�6�B� [�ޯ6�TŘ̓$�Ѭ|�oU=A�c	wk�C�2��{�
��lO�)l�#����g�i3Z��g�1O���@�ߤe�������(x�/o�*�V�i嫘uPz���pC����H�Ҁ�2�MY���I�@�_Il΅Eb��\\��i=v�ؒ9�����!1,B�����ߠc�����;��y>ވ Eo,1	ٓ2�u�1��u�G������� �2|��D��蓋lM��s,��obϸ��t³�X`̽�����,�G��)
��*�5h�r�3��XT���FL`W����
���#1����vF>���hnb�^R]}="�QÊ�Y�@��>��$��l�����S�ZM��*�,����=��ЊO�z?���G0����5����?�"A]��B�<��s�qwT�'� _ۥD��EJa�G-L�a��O�o#��
�[��t��V)!p���V�z> 2YF"�}�д�$���&�����/�2�ݖf���_~V�T"��	������ؖ�)����1-�������*�q<fZ�,�f�
�XsL���흎�Br����b<a����i�d���ґ��C
��'�neh%�|k^��
�|	Tڂ
�XY�(%`j9%��/�y�,' FT���]�3)_��f��T����
�Y���@Xv$��Wc�����3��Gǣy��䗸��j�����q�fWXt\t}�������kp[Q�S�W.�����*�C���D�J���p
�=�J噏$#}��]Ջ�əZv�� �~�Ԫ83*v�v:~؂#����L�8��x�sm�J' �Ё�a����� �N��,�a�j{z ��C��e0\@��V}&�"ь�����`�p��=�i���8x/l��W��_�)���2�p��<5g��7�$�%��Z�PP�)��@�3����Є�W��(�� p� ;� ��/���  4`����0�<�I!�۠��?�R��_��� 6        1Q !@A0Pa���q��"2�BRb�`������ 	? �E�!�J65��",<�TE��*�Ϙ�QP)�1�8	��cT�l,�E�"�#ppf�E����d�<!a
8'FzTBًP�|����P�!�h@g�p/�TOTJ+eC:=���0���܂1�g�E�s��! ���Q獡{'F{��T��T,0G6l�	@��	��'G��kG7
u���Q*( s��,	�:�80�UG���aEQEQE�D"�B!pX2��EQEQ�vy��{�\�p�p�p�p��&�	�{��4��&��)���M=�P60�MpA���РG��by-�
�&Ay�4 �
���.bt�/�����^̑B#�P�:����!}�X�� w��A)�4&�&�B {#wشH� w��}��mz)o����1�7Rv�A�}f�i�@Ј������㸭�7=�m����k�{Q��OoTDL�$@&A�I
�Eo�rߍ�QZF��}0v��^�g�I_E���*�M�#�~G� �s��E���E�鐕��(M8��꾣�(`�0�+�qَ>�_al�,ǲn�\ߛ�oTD+��c+޶Q�� �'���q&N�y�
�X`�n���	�ѫ�}�;���
?�]�B�S\]���X��Tz�� �?y�G�R����1���&$��BZ'D�憈�G�ql������y،v9���[#� H�8��u���6�Gk��_�"�_�]�;.~%��E����#��@7����GT����'l� D�:.杲5�8�#�t��Q0��d14Xc,��W!:#�<��W#������Gg�c�u��
i��!��-.�ި�B!d!�b��5���)����V���Gg�lMSB:� �SZ�;��� )���`��;���� 7�m'�{�X�+0:�N��32��Ի�d|�}���vjz����^b����{g�OS�����|�d���;��֦��k{����h��M	�4&�4&�ЀM	�4&��ܞ	�x7�~�5�5���S�V�3U�[��V�ru����']�oW#[+���ަ�W{\�l���������������� 0        !1@Q 0PAa2q"`��b������� 	? ��1�F�pE~�%��
��7�Ê'�/%�E�B(���A�EQ�:'���EOpB���(h%�p�����^K�G�r�(�J<U�e��<)(��N��"�P(
�QQy���@&S)��	��	� �o�v7�CYU9ߘ�|��_��/�J��5]�ޖ;�)����.g�"j�mV�Z�P1�d�`*� U����@��񱍼��VU _�T�_�PW��USU^�{�b�&�k��mb0]�<&}]���EΊX	�/��U.Y(� eW2Uq�%���Jh�n U�A"�MQU�_+)��U��"	����R��z�ko�Rx�z�@D! ��fWz��C]��dPyL��W�A����Ƞ��?
��:�+�D��=A� ?R�Q������&��5)�Ne��ts�M����Ŝ��,$?;�RtTyZ?��`m+ۀ���U}xJ��SM&�M5�� ���	��)��)��)��(�Ji4�E�Q��Q;��N����b�@@kYCHj���:�ݞ�_�v�c`]�68���5cwy���.q���n������.q��X�ά;�Ջ;��ñ��|;��ά;&���� F�9?��PK   u��T�i��T  o     jsons/user_defined.json��oK�0ƿ���Z��Yھ2�!s� C�6��.�I�1F����9����=��s��5������ׂ�B�MЖk#��v�K b��JJ^�Üml��9k�Z�=(���/�j�D�)�q�1�̟:AS'Ɯ94#�`Y��2 ��r*M����Snr-�wv6� ����zu��3Y*��l7�0u��7���P�^�y�:�jgSq=Jø'��h��h�����rmgf�k�^T!�ȍiD��>���D�k��)ŧF+�q�����'��'�d��A���쀌d/�/��=�|y��t���y����q����	[�AH���F?�]�\ɑk׭�OPK
   u��T��ఒ  �#                   cirkitFile.jsonPK
   ���T�߳�  /             �  images/6130fba0-ab36-4597-90ea-7b17dabf0cf4.jpgPK
   u��T�i��T  o               � jsons/user_defined.jsonPK      �   5   